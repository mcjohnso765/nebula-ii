* NGSPICE file created from team_01.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt team_01 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_out[0] gpio_out[10] gpio_out[11]
+ gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18]
+ gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24]
+ gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30]
+ gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6]
+ gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ _04789_ _04950_ _04951_ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or4_1
X_06883_ net962 cpu.RF0.registers\[2\]\[27\] net770 vssd1 vssd1 vccd1 vccd1 _02174_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11834__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ net1107 cpu.RF0.registers\[18\]\[3\] net853 vssd1 vssd1 vccd1 vccd1 _03913_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13840__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08553_ net1105 cpu.RF0.registers\[18\]\[5\] net853 vssd1 vssd1 vccd1 vccd1 _03844_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout162_A _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__inv_2
XANTENNA__07298__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__B1 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ net1106 cpu.RF0.registers\[24\]\[7\] net871 vssd1 vssd1 vccd1 vccd1 _03775_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07837__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A1 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07435_ net977 cpu.RF0.registers\[1\]\[1\] net807 vssd1 vssd1 vccd1 vccd1 _02726_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout427_A _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ net977 cpu.RF0.registers\[6\]\[2\] net802 vssd1 vssd1 vccd1 vccd1 _02657_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07986__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _04391_ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08262__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07297_ cpu.RF0.registers\[19\]\[4\] net615 net595 cpu.RF0.registers\[7\]\[4\] _02585_
+ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a221o_1
XANTENNA__14346__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13220__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1336_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ net952 cpu.RF0.registers\[12\]\[31\] net765 vssd1 vssd1 vccd1 vccd1 _04327_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07470__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 cpu.RF0.registers\[19\]\[8\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__A1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 cpu.RF0.registers\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 cpu.RF0.registers\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold373 cpu.RF0.registers\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_X clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 cpu.RF0.registers\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13370__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14496__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 cpu.RF0.registers\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net822 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
XANTENNA__08970__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout831 _02126_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_4
XANTENNA__12938__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ net625 _04863_ net1022 vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_70_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07507__B net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_4
Xfanout864 _02021_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
Xfanout875 _02010_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_8
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_4
X_09869_ _01785_ net717 net134 net632 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a31o_1
XANTENNA__07226__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1040 cpu.LCD0.row_2\[102\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 cpu.LCD0.row_1\[8\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11744__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_X clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1062 cpu.RF0.registers\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net2170 net247 net323 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
X_12880_ clknet_leaf_0_clk cpu.c0.next_count\[11\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[11\] sky130_fd_sc_hd__dfrtp_1
Xhold1073 cpu.RF0.registers\[16\]\[14\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 cpu.RF0.registers\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 cpu.RF0.registers\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ net2168 net236 net332 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__mux2_1
XANTENNA__14580__RESET_B net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__A1 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14550_ clknet_leaf_45_clk _01652_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[61\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07289__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ net1563 net138 net342 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08057__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13501_ clknet_leaf_89_clk _00614_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ cpu.LCD0.row_1\[119\] net1580 net905 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XANTENNA__10832__A1 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ clknet_leaf_30_clk cpu.RU0.next_write_i net1209 vssd1 vssd1 vccd1 vccd1 a1.WRITE_I
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ net1599 net149 net351 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ clknet_leaf_7_clk _00545_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ net2216 cpu.LCD0.row_1\[58\] net902 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08789__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ cpu.f0.write_data\[0\] _02716_ net995 vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__mux2_1
XANTENNA__09169__B _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__A0 cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ clknet_leaf_69_clk _00476_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12314_ cpu.LCD0.cnt_20ms\[1\] cpu.LCD0.cnt_20ms\[0\] net2922 vssd1 vssd1 vccd1 vccd1
+ _06196_ sky130_fd_sc_hd__a21o_1
XANTENNA__10060__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ clknet_leaf_33_clk cpu.RU0.next_FetchedData\[1\] net1248 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13713__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11919__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ cpu.LCD0.row_2\[69\] _05988_ _06015_ cpu.LCD0.row_1\[5\] vssd1 vssd1 vccd1
+ vccd1 _06141_ sky130_fd_sc_hd__a22o_1
XANTENNA__08005__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09202__A1 _03233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09202__B2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__A _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ cpu.LCD0.nextState\[5\] cpu.LCD0.nextState\[4\] cpu.LCD0.nextState\[3\] cpu.LCD0.nextState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__or4b_1
XFILLER_0_43_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08520__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11127_ net2256 net179 net421 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13863__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11058_ net2012 net164 net426 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08713__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net626 _05086_ net1023 vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09632__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14219__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11076__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14679_ net1401 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__08492__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13243__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14369__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07220_ net1034 cpu.RF0.registers\[31\]\[9\] net825 vssd1 vssd1 vccd1 vccd1 _02511_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07151_ net1043 cpu.RF0.registers\[17\]\[11\] net805 vssd1 vssd1 vccd1 vccd1 _02442_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10587__B1 _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07082_ cpu.RF0.registers\[19\]\[18\] net615 _02353_ _02355_ _02357_ vssd1 vssd1
+ vccd1 vccd1 _02373_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13393__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11829__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11000__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout127 _05148_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_2
XANTENNA__08952__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout149 net151 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
X_07984_ net1094 cpu.RF0.registers\[17\]\[28\] net884 vssd1 vssd1 vccd1 vccd1 _03275_
+ sky130_fd_sc_hd__and3_1
X_09723_ net486 _04798_ _04857_ _04384_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a221o_1
X_06935_ net958 cpu.RF0.registers\[15\]\[26\] net826 vssd1 vssd1 vccd1 vccd1 _02226_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10969__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12500__A1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11564__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _02437_ net300 vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__nand2_1
X_06866_ net966 net817 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__and2_1
XANTENNA__06885__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08605_ cpu.RF0.registers\[30\]\[4\] _02053_ _03894_ _03895_ net667 vssd1 vssd1 vccd1
+ vccd1 _03896_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08180__B2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12957__Q a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ net301 _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nor2_1
X_06797_ cpu.RF0.registers\[0\]\[30\] net661 net547 vssd1 vssd1 vccd1 vccd1 _02088_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__B1 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ cpu.RF0.registers\[4\]\[6\] net678 net639 cpu.RF0.registers\[26\]\[6\] _03813_
+ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12395__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ cpu.RF0.registers\[10\]\[8\] net692 _03755_ _03756_ _03757_ vssd1 vssd1 vccd1
+ vccd1 _03758_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07418_ net971 cpu.RF0.registers\[4\]\[0\] net783 vssd1 vssd1 vccd1 vccd1 _02709_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08398_ cpu.RF0.registers\[13\]\[10\] net657 net655 cpu.RF0.registers\[2\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08174__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire517 _02578_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_1
XANTENNA__13736__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07349_ _02631_ _02632_ _02638_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__or4_1
XANTENNA__08235__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10209__A cpu.IM0.address_IM\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1241_X net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1339_X net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ cpu.f0.i\[27\] cpu.f0.i\[28\] _05582_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10042__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09983__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11739__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09019_ cpu.RF0.registers\[10\]\[31\] net691 _04298_ _04299_ _04301_ vssd1 vssd1
+ vccd1 vccd1 _04310_ sky130_fd_sc_hd__a2111o_1
X_10291_ cpu.f0.i\[17\] _05526_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_72_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12424__A cpu.DM0.data_i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12030_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__inv_2
Xhold170 cpu.RF0.registers\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 cpu.RF0.registers\[4\]\[10\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 cpu.RF0.registers\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10750__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 _02058_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_8
Xfanout661 _02051_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout672 _02042_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_89_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09499__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout683 _02033_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_6
X_13981_ clknet_leaf_89_clk _01094_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout694 _02024_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_8
XANTENNA__11474__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12932_ clknet_leaf_29_clk _00121_ net1202 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10231__X _05484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__Q a1.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12863_ clknet_leaf_16_clk _00082_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13266__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14602_ clknet_leaf_52_clk _01704_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_11814_ net2603 net207 net334 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__mux2_1
X_12794_ net2895 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
X_14533_ clknet_leaf_48_clk _01635_ net1361 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[44\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10805__A1 cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11745_ net1648 net197 net342 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__mux2_1
XANTENNA__08474__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ clknet_leaf_22_clk _01574_ net1174 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ net2121 net212 net351 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ clknet_leaf_79_clk _00528_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08515__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10627_ net2528 net2365 net906 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__A _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ clknet_leaf_21_clk _01506_ net1176 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09908__A cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ clknet_leaf_11_clk _00459_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10558_ net1134 a1.ADR_I\[23\] net914 _05666_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ clknet_leaf_20_clk cpu.RU0.next_FetchedInstr\[16\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[16\] sky130_fd_sc_hd__dfrtp_1
X_10489_ net1494 net920 net749 a1.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 _00162_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07428__A cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12228_ cpu.LCD0.row_1\[108\] _06009_ _06031_ cpu.LCD0.row_1\[28\] _06124_ vssd1
+ vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10741__A0 cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ cpu.LCD0.row_2\[1\] _06016_ _06028_ cpu.LCD0.row_1\[113\] _06058_ vssd1 vssd1
+ vccd1 vccd1 _06059_ sky130_fd_sc_hd__a221o_1
XANTENNA__09643__A _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14041__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11384__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13609__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ net1096 net877 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06651_ a1.CPU_DAT_O\[19\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[19\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14191__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12246__B1 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06582_ cpu.LCD0.cnt_500hz\[9\] cpu.LCD0.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ _01957_ sky130_fd_sc_hd__and2_1
X_09370_ net305 _04657_ _04660_ _04648_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13759__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08321_ net942 cpu.RF0.registers\[6\]\[12\] net852 vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08252_ net1092 cpu.RF0.registers\[24\]\[15\] net871 vssd1 vssd1 vccd1 vccd1 _03543_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07203_ net969 cpu.RF0.registers\[1\]\[10\] net806 vssd1 vssd1 vccd1 vccd1 _02494_
+ sky130_fd_sc_hd__and3_1
X_08183_ net444 _03472_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout125_A _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__A cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07134_ cpu.RF0.registers\[4\]\[15\] net586 net566 cpu.RF0.registers\[11\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11559__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ net974 cpu.RF0.registers\[10\]\[18\] net788 vssd1 vssd1 vccd1 vccd1 _02356_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1034_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07728__A1 _03018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ cpu.RF0.registers\[11\]\[29\] net689 _03239_ _03244_ _03251_ vssd1 vssd1
+ vccd1 vccd1 _03258_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout661_A _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06896__B net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06951__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_A _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _04985_ _04991_ _04995_ _04996_ _04990_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__o2111a_1
X_06918_ _01850_ _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14172__RESET_B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08169__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ net1059 cpu.RF0.registers\[31\]\[29\] net828 net566 cpu.RF0.registers\[11\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_84_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07073__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__X _05131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ _02348_ net440 vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_65_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06849_ net963 cpu.RF0.registers\[3\]\[27\] net821 vssd1 vssd1 vccd1 vccd1 _02140_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12237__B1 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _04739_ _04858_ net482 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07801__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ net1105 cpu.RF0.registers\[28\]\[6\] net868 vssd1 vssd1 vccd1 vccd1 _03810_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ net277 _04784_ _04785_ _04788_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06467__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11530_ net2690 net143 net372 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08208__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ net2563 net157 net378 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XANTENNA__13311__Q cpu.DM0.data_i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ clknet_leaf_69_clk _00380_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10412_ cpu.f0.i\[18\] net268 vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14180_ clknet_leaf_96_clk _01293_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11392_ net2765 net153 net386 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11469__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10566__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ clknet_leaf_53_clk net2489 net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ cpu.f0.i\[24\] cpu.f0.i\[25\] _05567_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__and3_1
XANTENNA__10971__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10274_ net1417 _05520_ net726 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
X_13062_ clknet_leaf_54_clk _00242_ net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14064__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ cpu.RF0.registers\[30\]\[17\] net192 net310 vssd1 vssd1 vccd1 vccd1 _01417_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10723__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10402__A cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13964_ clknet_leaf_80_clk _01077_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08144__A1 cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ clknet_leaf_25_clk _00104_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10896__X _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13901__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07414__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ clknet_leaf_81_clk _01008_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08695__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11932__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12228__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ clknet_leaf_25_clk _00065_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08807__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09644__A1 _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08447__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ net1463 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ clknet_leaf_46_clk net2560 net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11728_ net2393 net140 net347 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14447_ clknet_leaf_25_clk _01557_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_11659_ net1574 net156 net354 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12400__B1 _06223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14378_ clknet_leaf_33_clk _01489_ net1247 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14407__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold906 _00314_ vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold917 cpu.RF0.registers\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13329_ clknet_leaf_74_clk _00442_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_38_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold928 cpu.RF0.registers\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__B1 _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 _01705_ vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10962__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ _02122_ _02946_ _02982_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__a21o_1
XANTENNA__13431__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14557__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ cpu.RF0.registers\[8\]\[22\] net611 _03083_ _03099_ _03100_ vssd1 vssd1 vccd1
+ vccd1 _03112_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10190__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net543 _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__or2_1
X_06703_ _01944_ _01949_ _01946_ cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 _00006_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__13581__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ cpu.RF0.registers\[8\]\[16\] net611 _02948_ _02967_ _02968_ vssd1 vssd1 vccd1
+ vccd1 _02974_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07324__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__S net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _04708_ _04712_ net485 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__mux2_1
XANTENNA__12219__B1 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ a1.CPU_DAT_O\[2\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[2\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07894__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__B cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07621__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _02275_ _03371_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__nand2_1
X_06565_ cpu.f0.read_i net987 _01948_ cpu.DM0.state\[2\] _01780_ vssd1 vssd1 vccd1
+ vccd1 _01949_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08438__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout242_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ _02832_ _02868_ net490 vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06496_ cpu.f0.state\[2\] _01875_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__and3_1
X_09284_ _03932_ _04496_ _04480_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ cpu.RF0.registers\[8\]\[14\] net707 net685 cpu.RF0.registers\[24\]\[14\]
+ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10982__A _03018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1249_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09938__A2 _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ net949 cpu.RF0.registers\[14\]\[20\] net840 vssd1 vssd1 vccd1 vccd1 _03457_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08452__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ cpu.RF0.registers\[0\]\[14\] net618 _02397_ _02407_ vssd1 vssd1 vccd1 vccd1
+ _02408_ sky130_fd_sc_hd__o22a_2
X_08097_ cpu.RF0.registers\[13\]\[22\] net659 net642 cpu.RF0.registers\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a22o_1
XANTENNA__09267__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload90 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload90/X sky130_fd_sc_hd__clkbuf_4
X_07048_ cpu.RF0.registers\[14\]\[19\] net576 _02329_ _02330_ _02331_ vssd1 vssd1
+ vccd1 vccd1 _02339_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07068__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1524_A a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10921__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08374__A1 _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__C_N _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10181__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13924__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ net448 _03269_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ net274 _05857_ _05858_ net926 net2581 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ net2446 cpu.LCD0.row_2\[94\] net1006 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XANTENNA__10484__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07885__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ clknet_leaf_74_clk _00793_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ _05332_ _05813_ net722 vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__mux2_2
XANTENNA__07090__X _02381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ net2392 net2173 net1005 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08429__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12562_ _01889_ _06313_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13235__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ clknet_leaf_66_clk _01414_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11513_ net2748 net210 net373 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__mux2_1
X_12493_ cpu.f0.i\[14\] _06277_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__or2_1
X_14232_ clknet_leaf_7_clk _01345_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11444_ net2619 net216 net378 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11199__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09177__B _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_68_clk _01276_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13454__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ net2505 net229 net387 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
X_13114_ clknet_leaf_55_clk _00294_ net1371 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ _05561_ _05564_ net307 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14094_ clknet_leaf_1_clk _01207_ net1142 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07409__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ clknet_leaf_51_clk _00225_ net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10257_ _01805_ _05500_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XANTENNA__10831__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1220 net1228 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07168__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07706__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10188_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nor2_1
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_2
Xfanout1264 net1265 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
Xfanout1275 net1300 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__clkbuf_4
Xfanout1286 net1287 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10132__A cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1297 net1299 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ clknet_leaf_92_clk _01060_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__A1 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09640__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_71_clk _00991_ net1341 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10786__B _05131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07441__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12829_ clknet_leaf_14_clk _00048_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[25\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12209__D _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08020_ net1097 cpu.RF0.registers\[18\]\[24\] net853 vssd1 vssd1 vccd1 vccd1 _03311_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold703 cpu.LCD0.row_2\[55\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 cpu.f0.num\[31\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 _00233_ vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 cpu.RF0.registers\[9\]\[0\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold747 cpu.RF0.registers\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 cpu.RF0.registers\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net717 net134 _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a21oi_1
Xhold769 cpu.RF0.registers\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07319__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13947__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload27_A clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ net1084 cpu.RF0.registers\[27\]\[27\] net880 vssd1 vssd1 vccd1 vccd1 _04213_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10741__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12152__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ cpu.RF0.registers\[2\]\[16\] net654 _04141_ _04142_ _04143_ vssd1 vssd1 vccd1
+ vccd1 _04144_ sky130_fd_sc_hd__a2111o_1
Xhold1403 cpu.RF0.registers\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 cpu.RF0.registers\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 cpu.LCD0.row_2\[11\] vssd1 vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06906__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1436 a1.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ net958 cpu.RF0.registers\[5\]\[22\] net796 vssd1 vssd1 vccd1 vccd1 _03095_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12971__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1447 cpu.RF0.registers\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ cpu.RF0.registers\[12\]\[18\] net697 _04058_ _04064_ _04068_ vssd1 vssd1
+ vccd1 vccd1 _04075_ sky130_fd_sc_hd__a2111o_1
Xhold1458 cpu.RF0.registers\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net2875 sky130_fd_sc_hd__dlygate4sd3_1
X_07735_ cpu.RF0.registers\[7\]\[20\] net595 _02167_ cpu.RF0.registers\[15\]\[20\]
+ _03023_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a221o_1
XANTENNA__08659__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11572__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ net1024 cpu.RF0.registers\[25\]\[16\] net756 vssd1 vssd1 vccd1 vccd1 _02957_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07989__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13327__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net292 _04409_ net305 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a21o_1
X_06617_ _01754_ _01753_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__nor2_1
X_07597_ net1046 cpu.RF0.registers\[24\]\[12\] net812 vssd1 vssd1 vccd1 vccd1 _02888_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1366_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__S net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ _04482_ _04626_ _04479_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a21o_1
X_06548_ _01780_ net1129 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08734__X _04025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08292__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _02311_ net445 vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__xnor2_1
X_06479_ cpu.K0.keyvalid _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__and2_2
XANTENNA__13477__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ _03507_ _03508_ net443 vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__a21boi_1
X_09198_ _04485_ _04488_ net484 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08613__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__inv_2
XANTENNA__08044__B1 _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10926__A0 cpu.DM0.readdata\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11160_ net2913 net152 net414 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07229__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11747__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ cpu.IM0.address_IM\[23\] _02310_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__or2_1
X_11091_ net1846 _05822_ net425 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12143__A2 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ net715 net132 _05316_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_41_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10154__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 cpu.DM0.readdata\[9\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 _01473_ vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net73 vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14102__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold63 net103 vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold74 _00180_ vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 cpu.LCD0.row_2\[121\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 net77 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_105_clk _00914_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12578__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__Q cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net2210 net136 net314 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__mux2_1
XANTENNA__09847__B2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13732_ clknet_leaf_96_clk _00845_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10944_ net2899 net927 _05682_ net275 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a22o_1
X_13663_ clknet_leaf_0_clk _00776_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875_ net723 _05273_ _05800_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ net2194 cpu.LCD0.row_2\[8\] net1008 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
XANTENNA__12603__A0 cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ clknet_leaf_93_clk _00707_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ cpu.K0.code\[4\] cpu.K0.code\[7\] cpu.K0.code\[6\] cpu.K0.code\[5\] vssd1
+ vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__or4b_2
XFILLER_0_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12476_ net262 _06266_ _06268_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__and3_1
XANTENNA__08092__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12844__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ clknet_leaf_78_clk _01328_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08523__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _05780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ net2869 net159 net383 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07389__A2 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ clknet_leaf_94_clk _01259_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11358_ net1824 net165 net390 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XANTENNA__11657__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__inv_2
XANTENNA__12994__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ clknet_leaf_87_clk _01190_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09635__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289_ net1942 net170 net398 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__mux2_1
XANTENNA__08338__A1 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__A2 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ clknet_leaf_54_clk _00000_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08889__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 net1053 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1062 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_2
Xfanout1083 net1085 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1094 net1109 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09838__A1 _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11392__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07520_ net1058 cpu.RF0.registers\[21\]\[6\] net797 vssd1 vssd1 vccd1 vccd1 _02811_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ net1055 cpu.RF0.registers\[17\]\[1\] net807 vssd1 vssd1 vccd1 vccd1 _02742_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06402_ net2827 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07382_ cpu.RF0.registers\[29\]\[2\] net601 _02655_ _02664_ _02667_ vssd1 vssd1 vccd1
+ vccd1 _02673_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09066__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ net484 _04409_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09052_ net952 cpu.RF0.registers\[4\]\[31\] net780 vssd1 vssd1 vccd1 vccd1 _04343_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_26_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12236__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ _03290_ _03291_ _03292_ _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__nor4_1
XFILLER_0_41_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold500 cpu.RF0.registers\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 cpu.RF0.registers\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10037__A cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 cpu.RF0.registers\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 cpu.RF0.registers\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold544 cpu.RF0.registers\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 cpu.RF0.registers\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold566 cpu.RF0.registers\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11567__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold577 cpu.RF0.registers\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold588 cpu.RF0.registers\[4\]\[18\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _05225_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__nor2_1
XANTENNA__14125__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold599 cpu.RF0.registers\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09526__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1114_A cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__A2 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13998__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ net490 _03019_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09885_ _05163_ _05165_ _05162_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a21o_1
Xhold1200 cpu.RF0.registers\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10136__B2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 cpu.LCD0.row_1\[24\] vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ net440 _04125_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__xor2_1
Xhold1222 cpu.RF0.registers\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 cpu.RF0.registers\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12832__SET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1244 cpu.RF0.registers\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 _00315_ vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 a1.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14275__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1277 cpu.RF0.registers\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net948 cpu.RF0.registers\[5\]\[18\] _02019_ vssd1 vssd1 vccd1 vccd1 _04058_
+ sky130_fd_sc_hd__and3_1
Xhold1288 cpu.RF0.registers\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1299 cpu.LCD0.row_1\[57\] vssd1 vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07718_ cpu.RF0.registers\[7\]\[17\] net596 _02986_ _02987_ _02995_ vssd1 vssd1 vccd1
+ vccd1 _03009_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ net668 _03972_ _03975_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07304__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07649_ net522 _02938_ _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o21ai_4
XANTENNA__10994__X _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07512__C net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ net1805 cpu.LCD0.row_1\[74\] net902 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09057__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ net296 net293 _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__mux2_1
XANTENNA__08265__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ net988 cpu.f0.write_data\[7\] vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__nor2_2
XANTENNA__08804__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__A3 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12809__RESET_B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ cpu.LCD0.cnt_20ms\[9\] _06203_ net1340 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07020__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ cpu.LCD0.row_1\[70\] _06001_ _06012_ cpu.LCD0.row_2\[110\] _06155_ vssd1
+ vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__a221o_1
X_14000_ clknet_leaf_74_clk _01113_ net1334 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11212_ net2596 net217 net406 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
X_12192_ _01773_ net743 _05989_ _06006_ cpu.LCD0.row_1\[35\] vssd1 vssd1 vccd1 vccd1
+ _06090_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11477__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
X_11143_ net2272 net229 net415 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XANTENNA__09455__B _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__A2 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__07256__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
X_11074_ net2740 net242 net423 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XANTENNA__14618__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10127__B2 cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10025_ _05278_ _05281_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_51_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09190__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13642__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ net2323 net198 net315 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08518__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ clknet_leaf_68_clk _00828_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ _05445_ _05838_ net721 vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__mux2_2
XANTENNA__07422__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11940__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13646_ clknet_leaf_5_clk _00759_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ cpu.DM0.readdata\[9\] _04846_ net736 vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__mux2_1
XANTENNA__08815__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13792__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ clknet_leaf_105_clk _00690_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_105_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ net2135 net560 net538 _05739_ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12528_ _06299_ _06300_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__nor2_1
XANTENNA__08253__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08008__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13022__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ cpu.f0.i\[2\] _06254_ net261 vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14148__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ clknet_leaf_77_clk _01242_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout309 _01936_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12107__A2 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07166__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ cpu.RF0.registers\[28\]\[26\] net578 _02228_ _02233_ _02235_ vssd1 vssd1
+ vccd1 vccd1 _02242_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14298__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _04840_ _04850_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__nand2b_1
X_06882_ net969 net771 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ net1101 cpu.RF0.registers\[20\]\[3\] net875 vssd1 vssd1 vccd1 vccd1 _03912_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net1106 cpu.RF0.registers\[25\]\[5\] net864 vssd1 vssd1 vccd1 vccd1 _03843_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07503_ net545 net510 _02761_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a21oi_4
XANTENNA__11135__B cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08495__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07332__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ net1106 cpu.RF0.registers\[23\]\[7\] net846 vssd1 vssd1 vccd1 vccd1 _03774_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11850__S net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07434_ net1055 cpu.RF0.registers\[22\]\[1\] net802 vssd1 vssd1 vccd1 vccd1 _02725_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__B net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07365_ net976 cpu.RF0.registers\[7\]\[2\] net819 vssd1 vssd1 vccd1 vccd1 _02656_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout322_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _02106_ _02115_ _02117_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09995__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07296_ cpu.RF0.registers\[8\]\[4\] net612 net584 cpu.RF0.registers\[2\]\[4\] _02586_
+ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a221o_1
XANTENNA__08163__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09035_ net1025 cpu.RF0.registers\[30\]\[31\] net761 vssd1 vssd1 vccd1 vccd1 _04326_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07470__A1 cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1231_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1329_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold330 cpu.RF0.registers\[18\]\[13\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 cpu.RF0.registers\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13515__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 cpu.RF0.registers\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 cpu.RF0.registers\[20\]\[0\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold374 cpu.RF0.registers\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 cpu.RF0.registers\[3\]\[26\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 cpu.RF0.registers\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07076__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ net127 _05221_ _05218_ net631 vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a211o_1
Xfanout832 net833 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09816__B1_N _05106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net856 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06981__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 _02019_ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
XANTENNA__13665__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _02004_ _05146_ _05157_ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__o211a_1
Xfanout898 net901 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_4
Xhold1030 cpu.RF0.registers\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1041 _01693_ vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _00232_ vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07804__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ cpu.RF0.registers\[1\]\[19\] net714 net650 cpu.RF0.registers\[14\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a22o_1
Xhold1063 cpu.RF0.registers\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _03045_ net444 net295 _05088_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a31o_1
Xhold1074 cpu.RF0.registers\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08178__Y _03469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 cpu.RF0.registers\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 cpu.LCD0.row_2\[50\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net505 _05910_ _05920_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and3_4
XFILLER_0_90_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07289__A1 cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net2873 net140 net343 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13314__Q cpu.DM0.data_i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13500_ clknet_leaf_11_clk _00613_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10712_ cpu.LCD0.row_1\[118\] net1642 net908 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XANTENNA__10293__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14480_ clknet_leaf_29_clk _00015_ net1209 vssd1 vssd1 vccd1 vccd1 cpu.RU0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11692_ net2663 net158 net350 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XANTENNA__10884__B net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13431_ clknet_leaf_65_clk _00544_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ net2743 net2705 net906 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__mux2_1
XANTENNA__08238__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13045__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ clknet_leaf_60_clk _00475_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10574_ net1135 net2368 net915 _05674_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ net1369 _05944_ _06195_ _05957_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_40_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ clknet_leaf_34_clk cpu.RU0.next_FetchedData\[0\] net1247 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07538__X _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ cpu.LCD0.row_2\[117\] _06007_ _06016_ cpu.LCD0.row_2\[5\] _06139_ vssd1 vssd1
+ vccd1 vccd1 _06140_ sky130_fd_sc_hd__a221o_1
XANTENNA__14440__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08801__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12175_ cpu.LCD0.row_2\[34\] _06004_ _06016_ cpu.LCD0.row_2\[2\] _06073_ vssd1 vssd1
+ vccd1 vccd1 _06074_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11126_ net2088 net154 net418 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07417__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__X _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06972__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11935__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ net1837 net169 net427 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14590__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ net126 _05286_ _05283_ net627 vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a211o_1
XANTENNA__10520__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11959_ net2763 net140 net320 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__mux2_1
XANTENNA__07152__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11670__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14678_ net1400 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_47_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08545__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06991__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13629_ clknet_leaf_90_clk _00742_ net1280 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08229__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09977__A0 cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07150_ net1050 cpu.RF0.registers\[30\]\[11\] net762 vssd1 vssd1 vccd1 vccd1 _02441_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10587__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13538__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__X _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07081_ cpu.RF0.registers\[27\]\[18\] net591 _02359_ _02364_ _02366_ vssd1 vssd1
+ vccd1 vccd1 _02372_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08280__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13688__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06512__B cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__A1 cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout128 net130 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
Xfanout139 _05843_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
X_07983_ net945 cpu.RF0.registers\[3\]\[28\] net836 vssd1 vssd1 vccd1 vccd1 _03274_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07327__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06963__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net301 _04909_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__nor2_1
X_06934_ net958 cpu.RF0.registers\[7\]\[26\] net816 vssd1 vssd1 vccd1 vccd1 _02225_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07183__X _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07624__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _04927_ _04943_ _04932_ _04934_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_2_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06865_ net963 cpu.RF0.registers\[13\]\[27\] net792 vssd1 vssd1 vccd1 vccd1 _02156_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout272_A _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ cpu.RF0.registers\[6\]\[4\] net675 _03872_ _03878_ _03879_ vssd1 vssd1 vccd1
+ vccd1 _03895_ sky130_fd_sc_hd__a2111o_1
X_09584_ net450 _04874_ _04873_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__o21a_1
XANTENNA__10050__A cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06796_ net1118 _02085_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__or2_2
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ cpu.RF0.registers\[9\]\[6\] net700 net658 cpu.RF0.registers\[13\]\[6\] _03817_
+ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a221o_1
XANTENNA__07062__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13068__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14313__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1279_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ net1095 cpu.RF0.registers\[31\]\[8\] net857 vssd1 vssd1 vccd1 vccd1 _03757_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07417_ net972 cpu.RF0.registers\[7\]\[0\] net818 vssd1 vssd1 vccd1 vccd1 _02708_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07691__A1 _02981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08397_ cpu.RF0.registers\[28\]\[10\] net705 net640 cpu.RF0.registers\[19\]\[10\]
+ _03687_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire507 _03795_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_1
Xwire518 _02575_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_1
X_07348_ cpu.RF0.registers\[5\]\[3\] _02148_ _02610_ _02611_ _02625_ vssd1 vssd1 vccd1
+ vccd1 _02639_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10578__A1 cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14463__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ cpu.RF0.registers\[27\]\[7\] net591 _02552_ _02559_ _02566_ vssd1 vssd1 vccd1
+ vccd1 _02570_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12905__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09018_ cpu.RF0.registers\[3\]\[31\] net642 _04296_ _04297_ _04305_ vssd1 vssd1 vccd1
+ vccd1 _04309_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07994__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ _01810_ _05527_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
XANTENNA__08190__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08621__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 cpu.FetchedInstr\[4\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 cpu.RF0.registers\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 cpu.RF0.registers\[31\]\[7\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 cpu.RF0.registers\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13309__Q cpu.DM0.data_i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout640 _02064_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 net653 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11755__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 _02051_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13980_ clknet_leaf_12_clk _01093_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 _02042_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09499__A2 _04784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 _02031_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_8
Xfanout695 _02024_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_4
X_12931_ clknet_leaf_29_clk _00120_ net1201 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12862_ clknet_leaf_16_clk _00081_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14601_ clknet_leaf_50_clk net2383 net1382 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_11813_ net1822 net174 net336 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__A1 _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12793_ net1553 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11490__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14532_ clknet_leaf_46_clk _01634_ net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12824__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11744_ net1652 net208 net345 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10805__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14463_ clknet_leaf_22_clk _01573_ net1174 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ cpu.RF0.registers\[20\]\[9\] net216 net350 vssd1 vssd1 vccd1 vccd1 _01089_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13414_ clknet_leaf_6_clk _00527_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net2226 cpu.LCD0.row_1\[40\] net909 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14394_ clknet_leaf_20_clk _01505_ net1176 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13345_ clknet_leaf_63_clk _00458_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10557_ net55 net919 vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10834__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08631__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09908__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07709__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13276_ clknet_leaf_16_clk cpu.RU0.next_FetchedInstr\[15\] net1196 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[15\] sky130_fd_sc_hd__dfrtp_1
X_10488_ net1518 net916 net751 a1.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12227_ cpu.LCD0.row_1\[36\] _06006_ _06037_ cpu.LCD0.row_1\[76\] vssd1 vssd1 vccd1
+ vccd1 _06124_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12191__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12158_ cpu.LCD0.row_2\[81\] _05990_ _06015_ cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1
+ vccd1 _06058_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06900__X _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10741__A1 _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13980__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net2711 net229 net420 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__mux2_1
XANTENNA__09643__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ net745 _05982_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__and3_4
XANTENNA_wire240_A _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06986__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13210__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ net2816 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06581_ _01955_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08320_ net1089 cpu.RF0.registers\[29\]\[12\] net849 vssd1 vssd1 vccd1 vccd1 _03611_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_50_clk_X clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13360__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12509__B cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ cpu.RF0.registers\[27\]\[15\] net712 net669 cpu.RF0.registers\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08870__B1 _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06507__B cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12928__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ cpu.RF0.registers\[3\]\[10\] net609 net583 cpu.RF0.registers\[6\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a22o_1
X_08182_ _02122_ _02946_ _03044_ _03121_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a211o_1
XANTENNA__10029__B cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07133_ net1050 cpu.RF0.registers\[31\]\[15\] net830 net583 cpu.RF0.registers\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a32o_1
XANTENNA__07425__A1 cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_X clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ net1063 cpu.RF0.registers\[28\]\[18\] net767 vssd1 vssd1 vccd1 vccd1 _02355_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1027_A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10732__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10732__B2 cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ cpu.RF0.registers\[5\]\[29\] net703 _03242_ _03246_ _03250_ vssd1 vssd1 vccd1
+ vccd1 _03257_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07354__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _04939_ _04940_ _04942_ _04921_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a31o_1
X_06917_ net741 _02004_ _02091_ net628 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__or4_4
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07897_ _03182_ _03184_ _03185_ _03187_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_84_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout654_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_84_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08153__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _04922_ _04925_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__or3_1
X_06848_ net966 net822 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_65_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ _04797_ _04857_ net471 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06779_ _02067_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout821_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout919_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net1106 cpu.RF0.registers\[30\]\[6\] net839 vssd1 vssd1 vccd1 vccd1 _03809_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_18_clk_X clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _04785_ _04786_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07113__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14141__RESET_B net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08616__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _03736_ _03737_ _03738_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or4_1
XANTENNA__08861__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07520__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13853__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ net1797 net162 net379 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ _01809_ net269 _05623_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_59_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11391_ net2449 net165 net386 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09810__C1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ clknet_leaf_56_clk _00310_ net1371 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07967__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ cpu.f0.i\[24\] _05567_ cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14209__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__A1 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08351__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14423__Q cpu.DM0.readdata\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ clknet_leaf_52_clk net2289 net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ net528 _05515_ _05516_ _05519_ net309 vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12173__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ net2929 net205 net310 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__mux2_1
XANTENNA__07719__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13039__Q cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13233__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14359__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 _02681_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout481 net483 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout492 _02121_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
X_13963_ clknet_leaf_90_clk _01076_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08144__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12914_ clknet_leaf_25_clk _00103_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13894_ clknet_leaf_5_clk _01007_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13383__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12845_ clknet_leaf_33_clk _00064_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ net2902 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07104__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ clknet_leaf_62_clk _01617_ net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11727_ net2308 net144 net348 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__mux2_1
XANTENNA__07430__C net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14446_ clknet_leaf_25_clk _01556_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_11658_ net2379 net161 net355 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10609_ net2178 cpu.LCD0.row_1\[23\] net904 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
X_14377_ clknet_leaf_33_clk _01488_ net1247 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09638__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11589_ net1798 net166 net362 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold907 cpu.RF0.registers\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 cpu.RF0.registers\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13328_ clknet_leaf_61_clk _00441_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_38_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold929 cpu.RF0.registers\[12\]\[30\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10962__A1 _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13259_ clknet_leaf_22_clk _00439_ net1172 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12164__B1 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10714__A1 a1.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11395__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07820_ cpu.RF0.registers\[7\]\[22\] net596 _03086_ _03091_ net621 vssd1 vssd1 vccd1
+ vccd1 _03111_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10190__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07751_ net1073 net633 net519 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a21o_2
XANTENNA_clkbuf_leaf_92_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
X_06702_ net34 net2627 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07682_ cpu.RF0.registers\[19\]\[16\] net616 _02954_ _02956_ _02964_ vssd1 vssd1
+ vccd1 vccd1 _02973_ sky130_fd_sc_hd__a2111o_1
X_09421_ _04709_ _04711_ net477 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__mux2_1
XANTENNA__12219__A1 cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06633_ a1.CPU_DAT_O\[1\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[1\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08717__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _03337_ _04641_ _03374_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__o21a_1
X_06564_ net987 _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08303_ net508 _03593_ cpu.IM0.address_IM\[13\] net551 vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__a2bb2o_4
X_09283_ net480 _04573_ _04481_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a21bo_1
X_06495_ _01880_ _01883_ _01884_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout235_A _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__A3 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ cpu.RF0.registers\[5\]\[14\] net703 net643 cpu.RF0.registers\[3\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10982__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ cpu.RF0.registers\[16\]\[20\] net637 _03453_ _03454_ _03455_ vssd1 vssd1
+ vccd1 vccd1 _03456_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout402_A _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07116_ _02402_ _02403_ _02404_ _02406_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08096_ cpu.RF0.registers\[27\]\[22\] net711 net699 cpu.RF0.registers\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a22o_1
XANTENNA__10953__A1 _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08171__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_12
XANTENNA_clkbuf_leaf_45_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload91/X sky130_fd_sc_hd__clkbuf_4
X_07047_ cpu.RF0.registers\[30\]\[19\] net565 _02322_ _02326_ _02332_ vssd1 vssd1
+ vccd1 vccd1 _02338_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_28_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1311_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14501__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _04287_ _04288_ _03304_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a21oi_2
X_07949_ net1097 cpu.RF0.registers\[29\]\[29\] net849 vssd1 vssd1 vccd1 vccd1 _03240_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14651__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07515__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_103_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ net986 cpu.f0.write_data\[10\] vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__or2_2
XANTENNA__08908__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _04909_ _04385_ net486 _04858_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ cpu.DM0.readdata\[18\] _05117_ net738 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12630_ net2146 cpu.LCD0.row_2\[24\] net1007 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08346__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ _06327_ net1639 _06320_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ net2487 net202 net372 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__mux2_1
X_14300_ clknet_leaf_15_clk _01413_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12492_ net263 _06276_ _06278_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__and3_1
XANTENNA__08643__A _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14031__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14231_ clknet_leaf_42_clk _01344_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11443_ cpu.RF0.registers\[13\]\[8\] net222 net379 vssd1 vssd1 vccd1 vccd1 _00864_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07259__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ clknet_leaf_60_clk _01275_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11374_ net2905 net232 net387 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ clknet_leaf_47_clk _00293_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[77\]
+ sky130_fd_sc_hd__dfstp_1
X_10325_ net1019 _05556_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__nor2_1
X_14093_ clknet_leaf_104_clk _01206_ net1156 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14181__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12146__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13044_ clknet_leaf_49_clk _00224_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ _05503_ _05504_ net309 vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or3b_1
XANTENNA__13749__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08365__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1221 net1223 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09193__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1268 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_2
X_10187_ _05448_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__o21ai_1
Xfanout1243 net1244 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07573__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
Xfanout1265 net1266 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12449__A1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1276 net1278 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__clkbuf_4
Xfanout1287 net1300 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_58_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10132__B _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11943__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1298 net1299 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_2
X_13946_ clknet_leaf_93_clk _01059_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14063__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09865__A2 _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13877_ clknet_leaf_73_clk _00990_ net1341 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09078__A0 _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12828_ clknet_leaf_42_clk _00047_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[24\]
+ sky130_fd_sc_hd__dfstp_4
XANTENNA__13129__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07160__C net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ net1430 net496 net281 cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09649__A _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ clknet_leaf_18_clk _01540_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13279__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14524__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 cpu.RF0.registers\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold715 cpu.RF0.registers\[20\]\[10\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold726 cpu.RF0.registers\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__A1 _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold737 cpu.RF0.registers\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _05250_ _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__xnor2_1
Xhold748 cpu.RF0.registers\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 cpu.RF0.registers\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ _04204_ _04211_ _03375_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12927__RESET_B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ net1074 cpu.RF0.registers\[31\]\[16\] net859 vssd1 vssd1 vccd1 vccd1 _04143_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12014__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06520__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1404 cpu.LCD0.row_2\[87\] vssd1 vssd1 vccd1 vccd1 net2810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 cpu.RF0.registers\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07564__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ net957 cpu.RF0.registers\[13\]\[22\] net791 vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__and3_1
Xhold1426 _01610_ vssd1 vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ _04071_ _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__or3_1
Xhold1437 cpu.RF0.registers\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net2843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1448 cpu.RF0.registers\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07335__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
Xhold1459 cpu.RF0.registers\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net2865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08108__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__S net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09305__B2 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ cpu.RF0.registers\[13\]\[20\] net598 net585 cpu.RF0.registers\[2\]\[20\]
+ _03024_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11112__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07632__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ net1025 cpu.RF0.registers\[27\]\[16\] net775 vssd1 vssd1 vccd1 vccd1 _02956_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ net292 _04409_ net306 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout1094_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06616_ _01984_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07596_ net1047 cpu.RF0.registers\[27\]\[12\] net776 vssd1 vssd1 vccd1 vccd1 _02887_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14054__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ net479 _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__nand2_1
XANTENNA__08166__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06547_ _01923_ _01935_ net1127 _01891_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__o211a_1
XANTENNA__12612__A1 cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07070__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ _03405_ _04555_ _03442_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a21o_1
XANTENNA__07095__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ _01867_ _01869_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08217_ _02945_ _03022_ _03044_ _03080_ net489 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__a311o_1
XFILLER_0_65_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09197_ net473 _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08044__A1 cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _03437_ _03438_ net445 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout986_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08079_ cpu.RF0.registers\[0\]\[25\] net664 net548 vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12128__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ cpu.IM0.address_IM\[22\] net930 _05379_ _05380_ vssd1 vssd1 vccd1 vccd1 _00045_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09294__A _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ net2504 net184 net423 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__B1_N net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _05298_ _05303_ _05315_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10233__A cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 _00170_ vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10154__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 _01525_ vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 net101 vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _00152_ vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 _00160_ vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 a1.CPU_DAT_I\[24\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold86 _01712_ vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_99_clk _00913_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 _00165_ vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ net2006 net142 net317 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07542__A cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ net1688 net927 _05680_ net275 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a22o_1
X_13731_ clknet_leaf_77_clk _00844_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ cpu.DM0.readdata\[13\] net736 net720 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__o21a_1
X_13662_ clknet_leaf_84_clk _00775_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06530__B2 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12613_ net2631 cpu.LCD0.row_2\[7\] net1002 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__mux2_1
XANTENNA__12594__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13593_ clknet_leaf_92_clk _00706_ net1240 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13421__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14547__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ _01888_ cpu.K0.code\[1\] cpu.K0.code\[0\] vssd1 vssd1 vccd1 vccd1 _06312_
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12475_ net1021 net257 vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__nand2_4
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10408__A cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ net2212 net177 net384 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
X_14214_ clknet_leaf_7_clk _01327_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_6 cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13571__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10917__B2 _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ clknet_leaf_66_clk _01258_ net1294 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11938__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10842__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net2647 net167 net390 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12119__B1 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ cpu.f0.i\[19\] cpu.f0.i\[20\] _05539_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and3_2
X_14076_ clknet_leaf_11_clk _01189_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net2790 net186 net400 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__mux2_1
X_13027_ clknet_leaf_27_clk net1130 net1184 vssd1 vssd1 vccd1 vccd1 a1.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08338__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ net1490 _05490_ net727 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__mux2_1
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
XANTENNA__07010__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1062 net1064 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07155__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_4
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11673__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_2
XANTENNA__08548__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06994__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ clknet_leaf_105_clk _01042_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ net978 cpu.RF0.registers\[2\]\[1\] net772 vssd1 vssd1 vccd1 vccd1 _02741_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06401_ cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__inv_2
X_07381_ cpu.RF0.registers\[3\]\[2\] net610 _02646_ _02660_ _02662_ vssd1 vssd1 vccd1
+ vccd1 _02672_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_57_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09120_ _02758_ _04375_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08283__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ net952 cpu.RF0.registers\[10\]\[31\] net786 vssd1 vssd1 vccd1 vccd1 _04342_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13914__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__A1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06824__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12009__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08002_ cpu.RF0.registers\[7\]\[28\] net652 _03277_ _03282_ _03283_ vssd1 vssd1 vccd1
+ vccd1 _03293_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09449__S1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 cpu.RF0.registers\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold512 a1.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 cpu.RF0.registers\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold534 cpu.RF0.registers\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 cpu.RF0.registers\[24\]\[30\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold556 cpu.RF0.registers\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold567 cpu.RF0.registers\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold578 cpu.RF0.registers\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09953_ _05224_ _02833_ cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__and3b_1
Xhold589 cpu.RF0.registers\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09526__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08904_ _02946_ _02982_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nor2_1
X_09884_ _05171_ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 cpu.LCD0.row_1\[81\] vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 cpu.RF0.registers\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net440 _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nand2_1
Xhold1223 cpu.RF0.registers\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07065__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1234 cpu.RF0.registers\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11583__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 cpu.RF0.registers\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 cpu.RF0.registers\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ net1095 cpu.RF0.registers\[30\]\[18\] net839 vssd1 vssd1 vccd1 vccd1 _04057_
+ sky130_fd_sc_hd__and3_1
Xhold1267 cpu.RF0.registers\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 cpu.LCD0.row_1\[102\] vssd1 vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 cpu.LCD0.row_1\[40\] vssd1 vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08458__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ cpu.RF0.registers\[5\]\[17\] net603 _02999_ _03002_ _03005_ vssd1 vssd1 vccd1
+ vccd1 _03008_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ cpu.RF0.registers\[2\]\[1\] net656 _03985_ _03986_ _03987_ vssd1 vssd1 vccd1
+ vccd1 _03988_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_36_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13444__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07648_ net543 _02904_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout901_A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ net968 cpu.RF0.registers\[2\]\[12\] net770 vssd1 vssd1 vccd1 vccd1 _02870_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10927__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__B _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09318_ _03119_ _03402_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__and2_1
X_10590_ _05683_ cpu.LCD0.row_1\[6\] net896 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
XANTENNA__08193__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13594__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09249_ _03195_ net434 net288 _04538_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__o22a_1
XANTENNA__10072__B2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ cpu.LCD0.row_1\[102\] _06024_ _06036_ cpu.LCD0.row_1\[22\] vssd1 vssd1 vccd1
+ vccd1 _06155_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11758__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ net1992 net223 net408 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XANTENNA__09765__A1 _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ cpu.LCD0.row_1\[107\] _06009_ _06037_ cpu.LCD0.row_1\[75\] _06088_ vssd1
+ vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__a221o_1
XANTENNA__07776__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
X_11142_ net1794 net232 net415 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11073_ net1708 net245 net423 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__12730__X _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _05276_ _05290_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__nand2_1
XANTENNA__07824__X _03115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07272__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ net1682 net210 net315 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__mux2_1
X_13714_ clknet_leaf_70_clk _00827_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10926_ cpu.DM0.readdata\[28\] _04716_ net739 vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12811__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13937__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13645_ clknet_leaf_101_clk _00758_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10857_ net1709 net221 net432 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ net287 _05737_ _05738_ net1014 cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1
+ vccd1 _05739_ sky130_fd_sc_hd__a32o_1
X_13576_ clknet_leaf_97_clk _00689_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ _01818_ _06298_ net260 vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12961__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ cpu.f0.i\[1\] cpu.f0.i\[2\] _06250_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11668__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11409_ net2511 net225 net384 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XANTENNA__12353__A cpu.K0.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09646__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ net1121 net1515 net530 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 _01515_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10366__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ clknet_leaf_74_clk _01241_ net1321 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13317__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ cpu.RF0.registers\[27\]\[26\] net591 _02218_ _02224_ _02229_ vssd1 vssd1
+ vccd1 vccd1 _02241_ sky130_fd_sc_hd__a2111o_1
X_14059_ clknet_leaf_90_clk _01172_ net1278 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11315__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07881__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ net1073 net1068 net1066 net1070 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_101_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13467__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ net1101 cpu.RF0.registers\[28\]\[3\] net869 vssd1 vssd1 vccd1 vccd1 _03911_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ net1105 cpu.RF0.registers\[24\]\[5\] net872 vssd1 vssd1 vccd1 vccd1 _03842_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_37_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07502_ _02789_ _02791_ _02792_ _02762_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__o31ai_2
XANTENNA__07298__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ net1106 cpu.RF0.registers\[30\]\[7\] net839 vssd1 vssd1 vccd1 vccd1 _03773_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12291__A2 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload87_A clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ net979 cpu.RF0.registers\[8\]\[1\] net813 vssd1 vssd1 vccd1 vccd1 _02724_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_18_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12087__X _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08725__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07364_ net1054 cpu.RF0.registers\[24\]\[2\] net813 vssd1 vssd1 vccd1 vccd1 _02655_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09103_ _04360_ net296 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09995__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07295_ cpu.RF0.registers\[29\]\[4\] net601 _02195_ cpu.RF0.registers\[30\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout315_A _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ net1025 cpu.RF0.registers\[29\]\[31\] net790 vssd1 vssd1 vccd1 vccd1 _04325_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07470__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__A _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09747__A1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11578__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 cpu.RF0.registers\[17\]\[28\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold331 cpu.RF0.registers\[22\]\[10\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1224_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 cpu.RF0.registers\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12751__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 cpu.RF0.registers\[20\]\[8\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 cpu.FetchedInstr\[6\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold375 cpu.RF0.registers\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14242__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 a1.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net814 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_4
Xhold397 cpu.RF0.registers\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08970__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__nor2_1
Xfanout822 net824 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10109__A2 _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout844 net847 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06981__A1 cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout855 _02035_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_4
Xfanout866 _02019_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
X_09867_ _05151_ _05156_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout851_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 cpu.RF0.registers\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_2
Xfanout899 net901 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
Xhold1031 cpu.RF0.registers\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 cpu.LCD0.row_2\[39\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 cpu.RF0.registers\[20\]\[2\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ cpu.RF0.registers\[21\]\[19\] net646 net645 cpu.RF0.registers\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a22o_1
XANTENNA__14392__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09798_ _03044_ net434 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08188__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1064 cpu.RF0.registers\[24\]\[18\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 cpu.RF0.registers\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 cpu.RF0.registers\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 cpu.RF0.registers\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ _03771_ _03801_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or3b_2
XANTENNA__07523__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11760_ net1734 net144 net343 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__mux2_1
XANTENNA__07289__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__X _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__A2 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ cpu.LCD0.row_1\[117\] cpu.LCD0.row_1\[125\] net899 vssd1 vssd1 vccd1 vccd1
+ _00341_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10657__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ net1665 net160 net351 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12438__A cpu.DM0.data_i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ net2555 net2370 net909 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux2_1
X_13430_ clknet_leaf_58_clk _00543_ net1368 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08354__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09986__A1 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_77_clk _00474_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08789__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ net64 net917 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07997__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ cpu.LCD0.cnt_20ms\[1\] cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _06195_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07461__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13292_ clknet_leaf_23_clk cpu.RU0.next_FetchedInstr\[31\] net1194 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[31\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06723__X _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11488__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ cpu.LCD0.row_2\[125\] _06022_ _06031_ cpu.LCD0.row_1\[29\] vssd1 vssd1 vccd1
+ vccd1 _06139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07267__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ cpu.LCD0.row_2\[26\] _06034_ _06036_ cpu.LCD0.row_1\[18\] vssd1 vssd1 vccd1
+ vccd1 _06073_ sky130_fd_sc_hd__a22o_1
XANTENNA__07213__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net1909 net165 net418 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ net2615 net182 net428 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _05284_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__nor2_1
XANTENNA__08713__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11958_ net1666 net147 net321 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07730__A _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10909_ cpu.DM0.readdata\[23\] _04577_ net734 vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__mux2_1
X_14677_ net1399 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__10823__A3 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ net2437 net159 net327 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__mux2_1
XANTENNA__14115__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13628_ clknet_leaf_12_clk _00741_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13559_ clknet_leaf_91_clk _00672_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ cpu.RF0.registers\[24\]\[18\] net607 net575 cpu.RF0.registers\[14\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14265__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11398__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10339__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07204__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout129 net130 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_2
X_07982_ net944 cpu.RF0.registers\[4\]\[28\] net875 vssd1 vssd1 vccd1 vccd1 _03273_
+ sky130_fd_sc_hd__and3_1
X_09721_ _04968_ _05011_ net272 _04712_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12857__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06933_ net958 cpu.RF0.registers\[3\]\[26\] net822 vssd1 vssd1 vccd1 vccd1 _02224_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09652_ _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__and2b_1
XANTENNA__12500__A3 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12022__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06864_ net983 net793 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08603_ cpu.RF0.registers\[1\]\[4\] net713 net686 cpu.RF0.registers\[31\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a22o_1
X_09583_ _04420_ _04431_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__or2_1
X_06795_ net1118 _02085_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__nor2_2
XANTENNA__10050__B _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ cpu.RF0.registers\[2\]\[6\] net656 _03822_ _03823_ _03824_ vssd1 vssd1 vccd1
+ vccd1 _03825_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_82_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12264__A2 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08465_ net946 cpu.RF0.registers\[14\]\[8\] net839 vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ net1048 cpu.RF0.registers\[26\]\[0\] net788 vssd1 vssd1 vccd1 vccd1 _02707_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ cpu.RF0.registers\[9\]\[10\] net701 net660 cpu.RF0.registers\[30\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire508 _03592_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14608__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ cpu.RF0.registers\[23\]\[3\] net613 _02612_ _02621_ net622 vssd1 vssd1 vccd1
+ vccd1 _02638_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1341_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07278_ cpu.RF0.registers\[16\]\[7\] net581 _02547_ _02554_ _02565_ vssd1 vssd1 vccd1
+ vccd1 _02569_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08640__A1 cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout899_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ cpu.RF0.registers\[8\]\[31\] net708 net640 cpu.RF0.registers\[19\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11101__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1227_X net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 a1.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 cpu.RF0.registers\[10\]\[30\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07518__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 cpu.LCD0.row_2\[123\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 cpu.DM0.readdata\[19\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 cpu.LCD0.row_1\[123\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10750__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout641 _02064_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_4
X_09919_ _05203_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__nor2_1
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_8
Xfanout663 net664 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout674 net676 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 _02031_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
X_12930_ clknet_leaf_29_clk _00119_ net1201 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout696 net698 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12861_ clknet_leaf_16_clk _00080_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13325__Q cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13012__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600_ clknet_leaf_52_clk net1898 net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14138__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11812_ net2116 net195 net336 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__mux2_1
XANTENNA__08646__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__X _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ net1418 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10266__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07550__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ clknet_leaf_61_clk net2456 net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11743_ net1842 net202 net343 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14462_ clknet_leaf_22_clk _01572_ net1179 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_12_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13162__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07682__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ net1759 net221 net353 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14288__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10018__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ clknet_leaf_8_clk _00526_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10625_ net2052 cpu.LCD0.row_1\[39\] net903 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__mux2_1
X_14393_ clknet_leaf_21_clk _01504_ net1176 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14088__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10556_ net1135 net2918 net915 _05665_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__a31o_1
X_13344_ clknet_leaf_8_clk _00457_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08381__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ net1469 net920 net749 a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__a22o_1
X_13275_ clknet_leaf_24_clk cpu.RU0.next_FetchedInstr\[14\] net1205 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11518__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12226_ _06116_ _06118_ _06120_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12157_ cpu.LCD0.row_1\[65\] _06001_ _06021_ cpu.LCD0.row_1\[89\] _06056_ vssd1 vssd1
+ vccd1 vccd1 _06057_ sky130_fd_sc_hd__a221o_1
XANTENNA__09483__Y _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10850__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11108_ net2510 net232 net420 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__mux2_1
X_12088_ cpu.LCD0.nextState\[1\] cpu.LCD0.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05989_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_21_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09344__C1 _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ net2467 net247 net429 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
XANTENNA__09895__B1 cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07163__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11681__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06580_ cpu.LCD0.cnt_500hz\[0\] cpu.LCD0.cnt_500hz\[1\] cpu.LCD0.cnt_500hz\[3\] cpu.LCD0.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__and4_1
XANTENNA__12246__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08556__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13505__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08250_ cpu.RF0.registers\[9\]\[15\] net700 net655 cpu.RF0.registers\[2\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08870__A1 _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10009__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07201_ net968 cpu.RF0.registers\[9\]\[10\] net757 vssd1 vssd1 vccd1 vccd1 _02492_
+ sky130_fd_sc_hd__and3_1
X_08181_ _02945_ _03022_ _03045_ net489 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13655__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ cpu.RF0.registers\[15\]\[15\] net590 net588 cpu.RF0.registers\[1\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07425__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06804__A cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07063_ net975 cpu.RF0.registers\[12\]\[18\] net767 vssd1 vssd1 vccd1 vccd1 _02354_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10422__C_N net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12017__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07338__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__S net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__Y _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _03243_ _03253_ _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__or4_1
XANTENNA__08138__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _04920_ _04989_ _04992_ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__o211a_1
XANTENNA__07354__B _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06916_ cpu.RF0.registers\[0\]\[27\] net617 _02203_ _02206_ vssd1 vssd1 vccd1 vccd1
+ _02207_ sky130_fd_sc_hd__o22a_4
XFILLER_0_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07896_ cpu.RF0.registers\[18\]\[29\] net579 net570 cpu.RF0.registers\[10\]\[29\]
+ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08169__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__B2 a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_4_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _03044_ net444 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__xnor2_1
X_06847_ net969 net813 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__and2_2
XANTENNA__07073__C net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12237__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _04822_ _04855_ net457 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__mux2_1
X_06778_ cpu.RF0.registers\[1\]\[30\] net714 net660 cpu.RF0.registers\[30\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__a22o_1
XANTENNA__13185__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ net1105 cpu.RF0.registers\[20\]\[6\] net875 vssd1 vssd1 vccd1 vccd1 _03808_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07801__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net298 _04786_ _04787_ _02473_ net291 vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08448_ cpu.RF0.registers\[20\]\[8\] net709 net695 cpu.RF0.registers\[17\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08379_ net1089 cpu.RF0.registers\[29\]\[10\] net850 vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14181__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ net1124 _01810_ net265 vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__or3_1
XANTENNA__14580__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11390_ net1935 net167 net389 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14110__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10341_ cpu.f0.i\[25\] _05571_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__and2_1
XANTENNA__10971__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ clknet_leaf_49_clk _00240_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ _05517_ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ net2687 net174 net312 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__mux2_1
XANTENNA__11766__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10670__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08129__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net464 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_4
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_8
X_13962_ clknet_leaf_102_clk _01075_ net1213 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_45_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13528__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ clknet_leaf_26_clk _00102_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ clknet_leaf_10_clk _01006_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12228__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ clknet_leaf_32_clk _00063_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08376__A _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__A1 _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08807__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07711__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ net2878 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ clknet_leaf_52_clk net2174 net1377 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11726_ net1628 net148 net346 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ clknet_leaf_25_clk _01555_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11657_ net1968 net177 net356 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_54_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10608_ net2336 cpu.LCD0.row_1\[22\] net908 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07407__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14376_ clknet_leaf_32_clk _01487_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12400__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11588_ net1768 net169 net363 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold908 cpu.RF0.registers\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ clknet_leaf_66_clk _00440_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10539_ net45 net919 vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__and2_1
Xhold919 cpu.RF0.registers\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10962__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__A cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ clknet_leaf_22_clk _00438_ net1171 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07158__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _05998_ _06000_ _06001_ _06004_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12361__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ clknet_leaf_36_clk _00369_ net1265 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14303__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06997__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07750_ cpu.RF0.registers\[0\]\[20\] net619 _03036_ _03040_ vssd1 vssd1 vccd1 vccd1
+ _03041_ sky130_fd_sc_hd__o22a_4
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06701_ cpu.LCD0.cnt_500hz\[13\] _01998_ cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1
+ vccd1 cpu.LCD0.lcd_en sky130_fd_sc_hd__a21oi_1
XANTENNA__14453__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ cpu.RF0.registers\[12\]\[16\] net572 _02950_ _02957_ _02958_ vssd1 vssd1
+ vccd1 vccd1 _02972_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06632_ a1.CPU_DAT_O\[0\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[0\]
+ sky130_fd_sc_hd__and2_1
X_09420_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__inv_2
XANTENNA__12219__A2 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__A2 _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06563_ cpu.DM0.enable _01779_ net736 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__or3_1
X_09351_ _03337_ _03374_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__nor3_1
XFILLER_0_74_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06518__B net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08302_ cpu.RF0.registers\[0\]\[13\] net662 net547 vssd1 vssd1 vccd1 vccd1 _03593_
+ sky130_fd_sc_hd__o21ai_1
X_09282_ _04571_ _04572_ net475 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__mux2_1
X_06494_ cpu.FetchedInstr\[12\] cpu.FetchedInstr\[15\] cpu.FetchedInstr\[14\] cpu.FetchedInstr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_72_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08573__X _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08233_ cpu.RF0.registers\[18\]\[14\] net681 net678 cpu.RF0.registers\[4\]\[14\]
+ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_A _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ net1099 cpu.RF0.registers\[18\]\[20\] net854 vssd1 vssd1 vccd1 vccd1 _03455_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07115_ cpu.RF0.registers\[16\]\[14\] net581 net573 cpu.RF0.registers\[9\]\[14\]
+ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a221o_1
XANTENNA__08452__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08095_ cpu.RF0.registers\[17\]\[22\] net694 _03378_ _03380_ _03381_ vssd1 vssd1
+ vccd1 vccd1 _03386_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08071__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload70/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__09845__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ cpu.RF0.registers\[24\]\[19\] net608 _02318_ _02325_ _02334_ vssd1 vssd1
+ vccd1 vccd1 _02337_ sky130_fd_sc_hd__a2111o_1
Xclkload81 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_2
Xclkload92 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__06821__X _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07068__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08359__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1304_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _04204_ _04211_ _04285_ _04286_ _03375_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_93_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07948_ net1098 cpu.RF0.registers\[19\]\[29\] net836 vssd1 vssd1 vccd1 vccd1 _03239_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout931_A _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ cpu.IG0.Instr\[28\] net634 _02210_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a21o_1
XANTENNA__08531__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_X net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ _04886_ _04908_ net457 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__mux2_1
XANTENNA__08196__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07885__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ net2770 net190 net430 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ _02544_ _03729_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12091__B1 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ net1128 cpu.DM0.data_i\[1\] _06307_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07637__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ net2043 net213 net372 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__mux2_1
XANTENNA__10665__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12491_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__inv_2
XANTENNA__06715__Y _02006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ clknet_leaf_70_clk _01343_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11442_ net2590 net226 net380 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14434__Q cpu.DM0.readdata\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14161_ clknet_leaf_77_clk _01274_ net1335 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11373_ net2543 net242 net387 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__mux2_1
XANTENNA__13200__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14326__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ clknet_leaf_49_clk _00292_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_10324_ _05560_ _05562_ net526 vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a21oi_1
X_14092_ clknet_leaf_68_clk _01205_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11496__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ clknet_leaf_45_clk _00223_ net1312 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10255_ cpu.f0.i\[12\] _05497_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nor2_1
XANTENNA__09474__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1200 net1210 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1386 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_4
XANTENNA__07022__B1 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13350__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14476__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_2
X_10186_ _05438_ _05440_ _05436_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a21oi_1
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07706__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1244 net1268 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
Xfanout1255 net1268 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08770__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12918__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1266 net1267 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_2
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_4
Xfanout290 _04407_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
Xfanout1288 net1291 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_4
Xfanout1299 net1300 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_2
X_13945_ clknet_leaf_13_clk _01058_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_64_clk_X clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload6_A clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07876__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ clknet_leaf_72_clk _00989_ net1340 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12827_ clknet_leaf_15_clk _00046_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09078__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ net1429 net496 net281 cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a22o_1
XANTENNA__08834__A _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_clk_X clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11709_ net1619 net213 net348 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XANTENNA__10575__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09649__B _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12689_ net2340 cpu.LCD0.row_2\[83\] net998 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
X_14428_ clknet_leaf_17_clk _01539_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12385__B2 cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold705 cpu.LCD0.row_1\[63\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14359_ clknet_leaf_71_clk _01472_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold716 cpu.RF0.registers\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 cpu.RF0.registers\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 cpu.RF0.registers\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 cpu.f0.num\[7\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
X_08920_ _03513_ _04210_ _04206_ _03440_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07185__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ net934 cpu.RF0.registers\[14\]\[16\] net837 vssd1 vssd1 vccd1 vccd1 _04142_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07616__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1405 cpu.RF0.registers\[11\]\[13\] vssd1 vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 cpu.RF0.registers\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ net958 cpu.RF0.registers\[14\]\[22\] net761 vssd1 vssd1 vccd1 vccd1 _03093_
+ sky130_fd_sc_hd__and3_1
Xhold1427 cpu.RF0.registers\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 cpu.RF0.registers\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13843__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ cpu.RF0.registers\[20\]\[18\] net710 net689 cpu.RF0.registers\[11\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a22o_1
Xhold1449 cpu.RF0.registers\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07913__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ net1055 cpu.RF0.registers\[31\]\[20\] net828 net602 cpu.RF0.registers\[5\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a32o_1
XANTENNA__08728__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ net1025 cpu.RF0.registers\[22\]\[16\] net799 vssd1 vssd1 vccd1 vccd1 _02955_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07867__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ net478 _04689_ _04691_ _04693_ net278 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10871__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13993__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06615_ net1350 _01972_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__nand2_1
X_07595_ net965 cpu.RF0.registers\[3\]\[12\] net821 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _04487_ _04624_ _04623_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a21oi_1
X_06546_ _01894_ _01901_ _01925_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06477_ cpu.K0.code\[2\] _01868_ cpu.K0.code\[3\] vssd1 vssd1 vccd1 vccd1 _01869_
+ sky130_fd_sc_hd__or3b_4
X_09265_ _03405_ _03442_ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout512_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13223__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14349__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _02122_ _02946_ _03079_ _03121_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__a2111o_1
X_09196_ net465 net437 _04486_ net453 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12376__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12376__B2 cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ net488 _03120_ _02312_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08044__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07647__X _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ net666 _03359_ _03364_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__or4_2
XANTENNA__14499__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13373__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout881_A _02008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout979_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ net1040 cpu.RF0.registers\[20\]\[19\] net781 vssd1 vssd1 vccd1 vccd1 _02320_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11169__X _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _05298_ _05303_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold10 cpu.f0.data_adr\[13\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07526__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 net120 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 net90 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _00158_ vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10801__X _05748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold54 cpu.f0.write_data\[31\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _00176_ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 cpu.RF0.registers\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 cpu.RF0.registers\[15\]\[0\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ net2125 net145 net316 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__mux2_1
XANTENNA__07542__B net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ clknet_leaf_95_clk _00843_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10942_ net1513 net927 _05678_ net275 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__a22o_1
XANTENNA__10311__B1 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A2 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14429__Q cpu.DM0.readdata\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ clknet_leaf_66_clk _00774_ net1282 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07261__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ net736 _04774_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__nand2_1
XANTENNA__06530__A2 cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__X _05932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ net2713 cpu.LCD0.row_2\[6\] net1006 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
X_13592_ clknet_leaf_19_clk _00705_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08654__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09102__X _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ _06309_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07491__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ net1021 net257 vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08092__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13716__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12367__B2 cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ clknet_leaf_9_clk _01326_ net1166 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ net2614 net154 net382 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08035__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13425__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14144_ clknet_leaf_9_clk _01257_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06461__X _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ net2537 net182 net391 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
XANTENNA__06902__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net1443 _05548_ net727 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
X_14075_ clknet_leaf_14_clk _01188_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13866__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11287_ net2305 net191 net398 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__mux2_1
X_13026_ clknet_leaf_29_clk _00215_ net1207 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
X_10238_ net307 _05485_ _05486_ _05489_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07436__C net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1030 net1033 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10143__B cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11954__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1044 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_2
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
X_10169_ net630 _04601_ net932 vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_2
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07292__X _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_1
XANTENNA__12890__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1096 net1109 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__buf_2
XFILLER_0_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13928_ clknet_leaf_99_clk _01041_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07849__A2 _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14213__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10853__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13859_ clknet_leaf_78_clk _00972_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06400_ cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ cpu.RF0.registers\[25\]\[2\] net568 _02649_ _02651_ _02652_ vssd1 vssd1 vccd1
+ vccd1 _02671_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_100_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ net952 cpu.RF0.registers\[2\]\[31\] net769 vssd1 vssd1 vccd1 vccd1 _04341_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10081__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12358__A1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ cpu.RF0.registers\[5\]\[28\] net703 net688 cpu.RF0.registers\[11\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a22o_1
XANTENNA__14641__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 cpu.c0.count\[15\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 cpu.RF0.registers\[13\]\[22\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07908__A cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 cpu.RF0.registers\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold535 cpu.RF0.registers\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload32_A clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 cpu.RF0.registers\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 cpu.RF0.registers\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _05233_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__or2_2
XANTENNA__12025__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold579 cpu.RF0.registers\[21\]\[3\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08903_ cpu.IM0.address_IM\[17\] net551 _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_
+ sky130_fd_sc_hd__a22o_4
X_09883_ cpu.IM0.address_IM\[4\] _02583_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout295_A _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08734__B1 _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 cpu.RF0.registers\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ _02348_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__xor2_2
Xhold1213 cpu.RF0.registers\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__A _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 cpu.RF0.registers\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 cpu.RF0.registers\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 cpu.FetchedInstr\[25\] vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 cpu.RF0.registers\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14021__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _03635_ _04049_ _04052_ _03567_ _04054_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1268 cpu.RF0.registers\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _00318_ vssd1 vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ net959 cpu.RF0.registers\[6\]\[17\] net799 vssd1 vssd1 vccd1 vccd1 _03007_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ cpu.RF0.registers\[30\]\[1\] _02053_ _02058_ cpu.RF0.registers\[14\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07647_ cpu.RF0.registers\[0\]\[13\] net620 _02933_ _02937_ vssd1 vssd1 vccd1 vccd1
+ _02938_ sky130_fd_sc_hd__o22a_2
XANTENNA__12548__X _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1371_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14171__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ cpu.CU0.funct3\[0\] _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13739__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ _03119_ _03402_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__nor2_1
X_06529_ cpu.f0.num\[8\] cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08265__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11104__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _03195_ net293 net448 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__or3b_1
XFILLER_0_84_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09179_ _04466_ _04469_ net457 vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__mux2_1
XANTENNA__13889__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11021__A1 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net2678 net227 net409 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
X_12190_ cpu.LCD0.row_1\[67\] _06001_ _06027_ cpu.LCD0.row_2\[43\] vssd1 vssd1 vccd1
+ vccd1 _06088_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ cpu.RF0.registers\[4\]\[4\] net241 net415 vssd1 vssd1 vccd1 vccd1 _00572_
+ sky130_fd_sc_hd__mux2_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__13119__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
X_11072_ net1757 net249 net423 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__07256__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13328__Q cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08649__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13269__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14514__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ net2029 net204 net315 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10835__A1 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ clknet_leaf_77_clk _00826_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08087__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ net2796 net148 net433 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13644_ clknet_leaf_74_clk _00757_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10856_ _05221_ _05787_ net721 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__mux2_2
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08384__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08815__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13575_ clknet_leaf_80_clk _00688_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08256__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10787_ net991 cpu.f0.data_adr\[21\] vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12526_ _01818_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__X _03962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__A_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ _06254_ _06255_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08008__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07216__A0 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11012__A1 _02247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ net1875 net228 net384 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
XANTENNA__06632__A a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ net1121 net2319 net530 cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14622__Q cpu.f0.write_data\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A1 cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__B2 cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ clknet_leaf_82_clk _01240_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ net2613 net248 net391 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XANTENNA__10771__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ clknet_leaf_100_clk _01171_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14044__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__A1 cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11684__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ clknet_leaf_34_clk _00198_ net1252 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06880_ net971 net783 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__and2_1
X_08550_ net1105 cpu.RF0.registers\[28\]\[5\] net869 vssd1 vssd1 vccd1 vccd1 _03841_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07750__X _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07501_ _02781_ _02782_ _02783_ _02784_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08481_ cpu.RF0.registers\[9\]\[7\] net700 net647 cpu.RF0.registers\[21\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a22o_1
XANTENNA__08495__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07432_ net1056 cpu.RF0.registers\[30\]\[1\] net764 vssd1 vssd1 vccd1 vccd1 _02723_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08725__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ net1054 cpu.RF0.registers\[26\]\[2\] net788 vssd1 vssd1 vccd1 vccd1 _02654_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10329__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ _02118_ _04391_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__A2 _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07294_ cpu.RF0.registers\[24\]\[4\] net607 net605 cpu.RF0.registers\[17\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ net952 cpu.RF0.registers\[6\]\[31\] net799 vssd1 vssd1 vccd1 vccd1 _04324_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11859__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__A1 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12200__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 cpu.RF0.registers\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 cpu.RF0.registers\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold332 cpu.RF0.registers\[14\]\[13\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 cpu.RF0.registers\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 cpu.RF0.registers\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__A0 cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 cpu.RF0.registers\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 a1.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold387 cpu.RF0.registers\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 cpu.RF0.registers\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _02145_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_8
X_09935_ cpu.IM0.address_IM\[8\] _05209_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__nor2_1
Xfanout812 net814 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_4
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
XANTENNA__07076__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10999__A _03115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08707__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08168__D1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_A _02037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net847 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
XANTENNA__06981__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14537__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ _05151_ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__nand2_1
XANTENNA__13411__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout867 net869 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_4
Xhold1010 cpu.LCD0.row_2\[17\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08469__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1021 cpu.RF0.registers\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _01951_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_1
X_08817_ _04095_ _04099_ _04103_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__or4_1
Xhold1032 cpu.RF0.registers\[13\]\[13\] vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 cpu.RF0.registers\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _03045_ net444 net296 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a21oi_1
Xhold1054 cpu.RF0.registers\[28\]\[16\] vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07804__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 cpu.LCD0.row_2\[73\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 cpu.RF0.registers\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _03870_ _04035_ _04036_ _03837_ _03803_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a311o_1
XFILLER_0_96_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1087 cpu.LCD0.row_1\[118\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 cpu.RF0.registers\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13561__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10817__A1 _04517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ net1103 cpu.RF0.registers\[23\]\[1\] net846 vssd1 vssd1 vccd1 vccd1 _03970_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_51_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ cpu.LCD0.row_1\[116\] cpu.LCD0.row_1\[124\] net904 vssd1 vssd1 vccd1 vccd1
+ _00340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06497__A1 cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11690_ net2350 net179 net352 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ net2441 net2333 net905 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__mux2_1
XANTENNA__08238__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__D cpu.RU0.next_read_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13360_ clknet_leaf_75_clk _00473_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10572_ net1135 net2939 net915 _05673_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__a31o_1
XANTENNA__09986__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08932__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11769__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ _01775_ net1369 _05957_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_40_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13291_ clknet_leaf_23_clk cpu.RU0.next_FetchedInstr\[30\] net1194 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[30\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12242_ cpu.LCD0.row_2\[109\] _06012_ _06133_ _06135_ _06137_ vssd1 vssd1 vccd1 vccd1
+ _06138_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09738__A2 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07548__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14067__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14442__Q cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ cpu.LCD0.row_2\[18\] _06003_ _06031_ cpu.LCD0.row_1\[26\] _06071_ vssd1 vssd1
+ vccd1 vccd1 _06072_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11124_ net1603 net169 net419 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13091__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06972__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ net2158 net172 net427 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10505__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08379__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ cpu.IM0.address_IM\[14\] _05271_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13904__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10520__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10848__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11957_ net2702 net150 net319 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10908_ net1558 net165 net433 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
X_14676_ net1398 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_47_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ net2707 net177 net328 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ clknet_leaf_14_clk _00740_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10839_ _05167_ _05775_ net721 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__mux2_4
XFILLER_0_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08229__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__A cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13558_ clknet_leaf_58_clk _00671_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08842__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11679__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ net1020 cpu.f0.i\[20\] _06286_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09657__B _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13489_ clknet_leaf_75_clk _00602_ net1334 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08937__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13434__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ net944 cpu.RF0.registers\[9\]\[28\] net863 vssd1 vssd1 vccd1 vccd1 _03272_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06963__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ net304 net436 net290 _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__o211a_1
XANTENNA__07464__Y _02755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06932_ net1029 cpu.RF0.registers\[23\]\[26\] net816 vssd1 vssd1 vccd1 vccd1 _02223_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07193__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13584__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _02312_ net445 _04922_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06863_ net1041 net787 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__and2_2
XANTENNA__07624__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ _03889_ _03890_ _03891_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12249__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ net455 _04421_ _04424_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__or3_1
X_06794_ _02082_ _02083_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__nand2_2
XFILLER_0_54_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08533_ cpu.RF0.registers\[3\]\[6\] net643 _03806_ _03808_ _03810_ vssd1 vssd1 vccd1
+ vccd1 _03824_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_82_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout160_A _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ net1095 cpu.RF0.registers\[16\]\[8\] net841 vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07415_ cpu.RF0.registers\[28\]\[0\] _02182_ _02704_ _02705_ net622 vssd1 vssd1 vccd1
+ vccd1 _02706_ sky130_fd_sc_hd__a2111o_1
X_08395_ net1089 cpu.RF0.registers\[16\]\[10\] net841 vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1167_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire509 _03230_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
X_07346_ _02633_ _02634_ _02635_ _02636_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07277_ net1060 cpu.RF0.registers\[24\]\[7\] net813 vssd1 vssd1 vccd1 vccd1 _02568_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1334_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08640__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10983__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09016_ cpu.RF0.registers\[24\]\[31\] net684 net654 cpu.RF0.registers\[2\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 cpu.DM0.readdata\[7\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _00159_ vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_X net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 cpu.RF0.registers\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _01714_ vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 cpu.f0.data_adr\[31\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _00339_ vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout620 _02128_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_4
Xfanout631 net632 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06954__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ cpu.IG0.Instr\[27\] cpu.IM0.address_IM\[7\] net520 vssd1 vssd1 vccd1 vccd1
+ _05204_ sky130_fd_sc_hd__and3_1
Xfanout642 net645 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout653 _02057_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _02051_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_6
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_8
X_09849_ net493 _05133_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a21oi_4
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12951__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ clknet_leaf_16_clk _00079_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08927__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13951__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ net2492 net198 net334 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12791_ net2529 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
X_14530_ clknet_leaf_51_clk _01632_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_11742_ net1737 net213 net343 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13307__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14437__Q cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14461_ clknet_leaf_23_clk _01571_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11673_ net2640 net226 net352 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ clknet_leaf_97_clk _00525_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ net2654 cpu.LCD0.row_1\[38\] net907 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XANTENNA__09758__A _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06734__X _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14392_ clknet_leaf_21_clk _01503_ net1180 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11499__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13343_ clknet_leaf_17_clk _00456_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_10555_ net54 net917 vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__and2_1
XANTENNA__13457__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08631__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13274_ clknet_leaf_24_clk cpu.RU0.next_FetchedInstr\[13\] net1204 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net102 net923 net748 net1556 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a22o_1
XANTENNA__07709__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ cpu.LCD0.row_1\[124\] _06014_ _06027_ cpu.LCD0.row_2\[44\] _06121_ vssd1
+ vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12191__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12156_ cpu.LCD0.row_1\[9\] _05994_ _06006_ cpu.LCD0.row_1\[33\] vssd1 vssd1 vccd1
+ vccd1 _06056_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11107_ net2749 net241 net420 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__mux2_1
XANTENNA__10432__A cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net746 _05982_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__and3_4
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11038_ net1959 net250 net429 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__mux2_1
XANTENNA__07444__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__A1 cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12989_ clknet_leaf_21_clk net1510 net1171 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13621__RESET_B net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07122__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14232__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14659_ net72 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ net1047 cpu.RF0.registers\[17\]\[10\] net805 vssd1 vssd1 vccd1 vccd1 _02491_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10009__A2 _05086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _03469_ _03470_ cpu.IM0.address_IM\[20\] net553 vssd1 vssd1 vccd1 vccd1 _03471_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07131_ _02412_ _02413_ _02414_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__or4_2
XFILLER_0_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14382__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06804__B cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07188__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ net1063 cpu.RF0.registers\[31\]\[18\] net829 vssd1 vssd1 vccd1 vccd1 _02353_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12182__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10193__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10732__A3 _05698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12974__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ cpu.RF0.registers\[28\]\[29\] net705 net646 cpu.RF0.registers\[21\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09703_ _04914_ _04993_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__nand2_1
X_06915_ _02197_ _02198_ _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ cpu.RF0.registers\[24\]\[29\] net607 net575 cpu.RF0.registers\[14\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a22o_1
XANTENNA__08689__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09634_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__inv_2
XANTENNA__10496__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06846_ net1073 net1071 net1068 net1066 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__nor4b_1
XANTENNA__06881__D_N net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07651__A _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09565_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06777_ cpu.RF0.registers\[18\]\[30\] net680 _02055_ _02015_ _02027_ vssd1 vssd1
+ vccd1 vccd1 _02068_ sky130_fd_sc_hd__a2111o_1
X_08516_ net1104 cpu.RF0.registers\[19\]\[6\] net836 vssd1 vssd1 vccd1 vccd1 _03807_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_61_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _03664_ net295 _04402_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07113__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08447_ cpu.RF0.registers\[27\]\[8\] net712 net672 cpu.RF0.registers\[29\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__a22o_1
XANTENNA__09849__Y _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08861__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout807_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _03664_ _03667_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08482__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08074__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ net1063 cpu.RF0.registers\[17\]\[3\] net806 vssd1 vssd1 vccd1 vccd1 _02620_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_59_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10956__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ cpu.f0.i\[25\] _05571_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ cpu.f0.i\[13\] cpu.f0.i\[14\] _05503_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__and3_1
XANTENNA__12173__A2 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07385__X _02676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net2022 net194 net312 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__mux2_1
XANTENNA__07826__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14105__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
Xfanout461 net464 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09326__B1 _04616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout472 _02681_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
X_13961_ clknet_leaf_2_clk _01074_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout483 _02643_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07264__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout494 _02119_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_4
XANTENNA__11782__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12912_ clknet_leaf_25_clk _00101_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07888__B1 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ clknet_leaf_98_clk _01005_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08657__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__A2 _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14255__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ clknet_leaf_31_clk _00062_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ net2830 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07104__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14513_ clknet_leaf_49_clk _01615_ net1376 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ net1800 net156 net346 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ clknet_leaf_27_clk _01554_ net1188 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_11656_ net2016 net154 net354 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12847__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10607_ cpu.LCD0.row_1\[13\] cpu.LCD0.row_1\[21\] net896 vssd1 vssd1 vccd1 vccd1
+ _00237_ sky130_fd_sc_hd__mux2_1
XANTENNA__08065__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375_ clknet_leaf_32_clk _01486_ net1250 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09801__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ net2638 net181 net365 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08604__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13326_ clknet_leaf_21_clk net892 net1177 vssd1 vssd1 vccd1 vccd1 cpu.DM0.ihit sky130_fd_sc_hd__dfrtp_1
X_10538_ net1134 net1913 net914 _05656_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__a31o_1
Xhold909 cpu.RF0.registers\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07439__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ clknet_leaf_43_clk _00437_ net1304 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12997__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ net19 net752 net562 net1858 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__o22a_1
XANTENNA__12164__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ cpu.LCD0.nextState\[3\] net743 _05989_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_
+ sky130_fd_sc_hd__a31o_1
X_13188_ clknet_leaf_36_clk _00368_ net1265 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06640__A a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ cpu.LCD0.row_1\[120\] _06014_ _06039_ net556 _06013_ vssd1 vssd1 vccd1 vccd1
+ _06040_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10162__A cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09951__A cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13873__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12321__C1 net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ cpu.LCD0.cnt_500hz\[8\] _01957_ _01997_ cpu.LCD0.cnt_500hz\[11\] cpu.LCD0.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a311o_1
XANTENNA__10478__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ cpu.RF0.registers\[10\]\[16\] net569 _02962_ _02965_ _02969_ vssd1 vssd1
+ vccd1 vccd1 _02971_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07879__B1 _02210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07343__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire510_A _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ _01971_ _01993_ _01995_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a21o_1
XANTENNA__13622__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ _04204_ _04211_ _03340_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a21oi_2
X_06562_ net1123 net988 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ _03582_ _03586_ _03590_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nor4_1
XFILLER_0_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09281_ net495 _03268_ net447 _04243_ net465 net454 vssd1 vssd1 vccd1 vccd1 _04572_
+ sky130_fd_sc_hd__mux4_1
X_06493_ cpu.FetchedInstr\[9\] cpu.FetchedInstr\[8\] cpu.FetchedInstr\[11\] cpu.FetchedInstr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__or4_1
XANTENNA__07500__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08232_ cpu.RF0.registers\[20\]\[14\] net709 net697 cpu.RF0.registers\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09829__C _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13772__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ net1099 cpu.RF0.registers\[21\]\[20\] net865 vssd1 vssd1 vccd1 vccd1 _03454_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09699__A_N net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07114_ cpu.RF0.registers\[5\]\[14\] net602 net599 cpu.RF0.registers\[26\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ net936 cpu.RF0.registers\[10\]\[22\] net860 vssd1 vssd1 vccd1 vccd1 _03385_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload60 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload60/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11867__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07045_ cpu.RF0.registers\[12\]\[19\] net572 _02327_ _02328_ _02333_ vssd1 vssd1
+ vccd1 vccd1 _02336_ sky130_fd_sc_hd__a2111o_1
Xclkload71 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload71/X sky130_fd_sc_hd__clkbuf_4
Xclkload82 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload82/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14128__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1032_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__12155__A2 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09020__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08996_ _04247_ _04282_ _04284_ _04279_ _04280_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__a311oi_4
XANTENNA__13152__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14278__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__inv_2
XANTENNA__12698__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10469__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ cpu.RF0.registers\[0\]\[28\] net619 _03159_ _03168_ vssd1 vssd1 vccd1 vccd1
+ _03169_ sky130_fd_sc_hd__o22ai_4
XANTENNA__10800__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__A _02865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _04465_ _04467_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__or2_1
X_06829_ _02112_ _02115_ _02117_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__or3_1
XANTENNA__07812__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _02544_ _03729_ net295 _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a31o_1
XANTENNA__08764__X _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09479_ net292 _04481_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or2_2
XFILLER_0_13_1427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ cpu.RF0.registers\[15\]\[9\] net216 net370 vssd1 vssd1 vccd1 vccd1 _00929_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ _05512_ _06264_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09101__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ net2329 net231 net380 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XANTENNA__10929__A0 cpu.DM0.readdata\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__A cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ clknet_leaf_75_clk _01273_ net1334 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11372_ net2658 net245 net387 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__mux2_1
XANTENNA__07259__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ clknet_leaf_46_clk net2254 net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11777__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ net540 _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__nand2_1
XANTENNA__07827__Y _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14091_ clknet_leaf_91_clk _01204_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12146__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ clknet_leaf_45_clk _00222_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07556__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ cpu.f0.i\[11\] cpu.f0.i\[12\] _05491_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1201 net1203 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1220 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_4
Xfanout1223 net1228 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
X_10185_ cpu.IM0.address_IM\[29\] _03193_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__and2_1
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
Xfanout1245 net1255 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net1267 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_4
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__clkbuf_4
Xfanout280 _01767_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout1278 net1283 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__clkbuf_4
Xfanout291 _04406_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
Xfanout1289 net1291 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13645__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ clknet_leaf_18_clk _01057_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13875_ clknet_leaf_67_clk _00988_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12826_ clknet_leaf_15_clk _00045_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13795__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10856__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12757_ cpu.f0.write_data\[15\] net499 net280 cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1
+ _01736_ sky130_fd_sc_hd__a22o_1
X_11708_ net1695 net216 net346 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
XANTENNA__06635__A a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12688_ net2374 cpu.LCD0.row_2\[82\] net1001 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08553__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09011__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14427_ clknet_leaf_18_clk _01538_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13025__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ net2626 net228 net356 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14358_ clknet_leaf_72_clk _01471_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 _00287_ vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 cpu.RF0.registers\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11687__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 cpu.f0.num\[19\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[16\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[16\] sky130_fd_sc_hd__dfrtp_1
X_14289_ clknet_leaf_76_clk _01402_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold739 cpu.RF0.registers\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__A2 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06370__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10148__B2 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14420__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08210__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net1074 cpu.RF0.registers\[27\]\[16\] net880 vssd1 vssd1 vccd1 vccd1 _04141_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08761__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1406 cpu.RF0.registers\[8\]\[29\] vssd1 vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
X_07801_ net957 cpu.RF0.registers\[10\]\[22\] net786 vssd1 vssd1 vccd1 vccd1 _03092_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07564__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1417 cpu.RF0.registers\[24\]\[1\] vssd1 vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ cpu.RF0.registers\[4\]\[18\] net678 _04059_ _04065_ _04069_ vssd1 vssd1 vccd1
+ vccd1 _04072_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1428 cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1439 cpu.RF0.registers\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
X_07732_ cpu.RF0.registers\[3\]\[20\] net610 net587 cpu.RF0.registers\[4\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_1
XANTENNA__14570__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06568__A_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08728__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ net953 cpu.RF0.registers\[11\]\[16\] net775 vssd1 vssd1 vccd1 vccd1 _02954_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07632__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06529__B cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ net449 _04509_ _04692_ _04384_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o211ai_1
X_06614_ _01970_ _01982_ _01983_ _01979_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a31o_1
X_07594_ net965 cpu.RF0.registers\[7\]\[12\] net817 vssd1 vssd1 vccd1 vccd1 _02885_
+ sky130_fd_sc_hd__and3_1
X_09333_ net474 _04483_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06545_ _01913_ _01930_ _01932_ _01933_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__or4b_1
XANTENNA__08816__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ _04205_ _04553_ _03407_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a21o_1
X_06476_ cpu.K0.code\[1\] cpu.K0.code\[0\] vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08215_ net488 _03044_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08029__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ net495 net460 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1247_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08146_ net488 _02312_ _03120_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or3_1
XANTENNA__13518__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09575__B _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ cpu.RF0.registers\[27\]\[25\] net711 _03365_ _03366_ _03367_ vssd1 vssd1
+ vccd1 vccd1 _03368_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_8_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12128__A2 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ net1040 cpu.RF0.registers\[22\]\[19\] net801 vssd1 vssd1 vccd1 vccd1 _02319_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10139__A1 cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07807__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__C net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13668__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 cpu.f0.data_adr\[16\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 cpu.RF0.registers\[0\]\[8\] vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 _00177_ vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 net96 vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ cpu.RF0.registers\[31\]\[26\] net687 net660 cpu.RF0.registers\[30\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 cpu.DM0.readdata\[12\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net76 vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net74 vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net1610 net150 net315 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__mux2_1
Xhold99 net85 vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10941_ net1782 net926 _05677_ net274 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13660_ clknet_leaf_8_clk _00773_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10862__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ net1888 net210 net430 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XANTENNA__08935__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12611_ cpu.LCD0.row_2\[13\] cpu.LCD0.row_2\[5\] net1000 vssd1 vssd1 vccd1 vccd1
+ _01604_ sky130_fd_sc_hd__mux2_1
XANTENNA__13048__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ clknet_leaf_64_clk _00704_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09465__C1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12542_ cpu.K0.code\[5\] cpu.K0.code\[7\] cpu.K0.code\[6\] cpu.K0.code\[4\] vssd1
+ vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__or4b_1
XANTENNA__06818__A1 cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12473_ net1021 _06264_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__or2_1
X_14212_ clknet_leaf_97_clk _01325_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13198__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ net2004 net165 net382 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06742__X _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14443__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_106_clk _01256_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11355_ net2665 net171 net393 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06902__B net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _05544_ _05546_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08991__A1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14074_ clknet_leaf_93_clk _01187_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11286_ net2783 net207 net398 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__mux2_1
X_13025_ clknet_leaf_29_clk _00214_ net1203 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13465__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10237_ _05487_ _05488_ net527 vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__and3b_1
XANTENNA__14593__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1020 cpu.f0.i\[19\] vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_2
XANTENNA__10143__C _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1031 net1033 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_2
XANTENNA__07573__X _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09940__B1 cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1044 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_2
Xfanout1053 net1064 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
X_10168_ net126 _05427_ _05433_ net630 vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1064 cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_1
Xfanout1086 net1091 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_2
X_10099_ cpu.IM0.address_IM\[22\] _03116_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09006__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08548__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ clknet_leaf_80_clk _01040_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07452__C net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11970__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13858_ clknet_leaf_95_clk _00971_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ clknet_leaf_37_clk _00028_ net1266 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08259__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13789_ clknet_leaf_67_clk _00902_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06365__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08000_ cpu.RF0.registers\[15\]\[28\] net683 net681 cpu.RF0.registers\[18\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a22o_1
XANTENNA__09759__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold503 cpu.RF0.registers\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07467__Y _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 cpu.RF0.registers\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07908__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold525 cpu.RF0.registers\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 cpu.RF0.registers\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 cpu.RF0.registers\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11210__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire842_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ cpu.CU0.bit30 cpu.IM0.address_IM\[10\] net520 vssd1 vssd1 vccd1 vccd1 _05234_
+ sky130_fd_sc_hd__and3_1
Xhold558 cpu.RF0.registers\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 cpu.RF0.registers\[6\]\[22\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload25_A clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ cpu.RF0.registers\[0\]\[17\] net661 net547 vssd1 vssd1 vccd1 vccd1 _04193_
+ sky130_fd_sc_hd__o21a_1
X_09882_ cpu.IM0.address_IM\[4\] _02583_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__and2_1
XANTENNA__08734__A1 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _02383_ _02945_ _03020_ net489 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__a31o_1
XANTENNA__07924__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1203 cpu.RF0.registers\[5\]\[26\] vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout190_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1214 cpu.RF0.registers\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 cpu.LCD0.row_2\[15\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13960__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1236 cpu.RF0.registers\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _03635_ _03801_ _04039_ _04047_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or4bb_4
XANTENNA__10350__A cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1247 cpu.RF0.registers\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 cpu.RF0.registers\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 cpu.RF0.registers\[4\]\[27\] vssd1 vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ net1027 cpu.RF0.registers\[27\]\[17\] net775 vssd1 vssd1 vccd1 vccd1 _03006_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08458__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__C net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ cpu.RF0.registers\[6\]\[1\] net675 net637 cpu.RF0.registers\[16\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11880__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14316__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07646_ _02928_ _02934_ _02935_ _02936_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06827__X _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07577_ _02473_ _02508_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ net485 _04488_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06528_ cpu.f0.num\[18\] _01811_ cpu.f0.num\[14\] _01806_ vssd1 vssd1 vccd1 vccd1
+ _01917_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14466__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1472_A cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09247_ _03196_ net448 vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nor2_1
X_06459_ cpu.RU0.state\[6\] net1130 a1.WRITE_I vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12908__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09178_ _04467_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout991_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ cpu.RF0.registers\[12\]\[23\] net696 net651 cpu.RF0.registers\[7\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a22o_1
XANTENNA__11021__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_X clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ net1915 net246 net415 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_11071_ net2884 net254 net424 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__07528__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_X clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ cpu.IM0.address_IM\[16\] _02947_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ net1700 net214 net316 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__mux2_1
XANTENNA__07272__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__A1 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13712_ clknet_leaf_74_clk _00825_ net1334 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10924_ _02001_ _05427_ _05835_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a22o_1
XANTENNA__06737__X _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ cpu.DM0.readdata\[8\] _04863_ net739 vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__mux2_1
X_13643_ clknet_leaf_86_clk _00756_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13574_ clknet_leaf_9_clk _00687_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ net991 _05131_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nand2_1
XANTENNA__08952__X _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12525_ cpu.f0.i\[26\] _06296_ _06298_ net260 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__o211a_1
XANTENNA__09767__Y _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13833__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ cpu.f0.i\[1\] _06250_ net263 vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_10_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07216__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ net2722 net235 net384 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11012__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ net1121 net1706 net530 cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 _01513_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06632__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14126_ clknet_leaf_2_clk _01239_ net1142 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12760__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ net1868 net250 net391 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10771__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__C net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10771__B2 cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ clknet_leaf_105_clk _01170_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ _05906_ net504 _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__and3_4
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13008_ clknet_leaf_34_clk _00197_ net1250 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09913__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14339__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13213__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07500_ net1061 cpu.RF0.registers\[31\]\[5\] net828 _02790_ net622 vssd1 vssd1 vccd1
+ vccd1 _02791_ sky130_fd_sc_hd__a311o_1
X_08480_ _03769_ _03770_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13363__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14489__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ net978 cpu.RF0.registers\[7\]\[1\] net818 vssd1 vssd1 vccd1 vccd1 _02722_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07910__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06807__B cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11205__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07362_ net1054 cpu.RF0.registers\[22\]\[2\] net803 vssd1 vssd1 vccd1 vccd1 _02653_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ _02118_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07293_ cpu.RF0.registers\[20\]\[4\] net594 net579 cpu.RF0.registers\[18\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
X_09032_ cpu.IM0.address_IM\[31\] net551 _04321_ _04322_ vssd1 vssd1 vccd1 vccd1 _04323_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 cpu.FetchedInstr\[29\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11003__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold311 cpu.RF0.registers\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 cpu.RF0.registers\[31\]\[10\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 cpu.RF0.registers\[17\]\[31\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__B1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12751__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold344 cpu.DM0.readdata\[30\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 cpu.RF0.registers\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07357__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold366 cpu.RF0.registers\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__A1 _05086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06966__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold377 cpu.RF0.registers\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold388 cpu.RF0.registers\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net803 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
X_09934_ cpu.IM0.address_IM\[8\] _05209_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__and2_2
Xhold399 cpu.LCD0.row_1\[66\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1112_A cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout824 _02131_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10999__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07654__A _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
X_09865_ cpu.IM0.address_IM\[0\] _02682_ _05154_ _05152_ vssd1 vssd1 vccd1 vccd1 _05156_
+ sky130_fd_sc_hd__a31o_1
Xfanout857 _02029_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_4
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 cpu.RF0.registers\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
Xhold1011 cpu.RF0.registers\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net881 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_8
Xhold1022 cpu.LCD0.row_1\[19\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 cpu.LCD0.row_2\[111\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ cpu.RF0.registers\[11\]\[19\] net690 _04104_ _04105_ _04106_ vssd1 vssd1
+ vccd1 vccd1 _04107_ sky130_fd_sc_hd__a2111o_1
X_09796_ _03477_ _04203_ _04210_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__nand3_1
Xhold1044 cpu.RF0.registers\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 cpu.LCD0.row_1\[10\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 _01664_ vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ _03870_ _04035_ _04036_ _03837_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__a31o_1
XANTENNA__12267__A1 cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 cpu.LCD0.row_2\[82\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13706__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1088 cpu.RF0.registers\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12559__X _06326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 cpu.RF0.registers\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ net1103 cpu.RF0.registers\[18\]\[1\] net853 vssd1 vssd1 vccd1 vccd1 _03969_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08485__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ net1045 cpu.RF0.registers\[19\]\[13\] net821 vssd1 vssd1 vccd1 vccd1 _02920_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_X net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13856__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10640_ net2185 net2937 net907 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__mux2_1
X_10571_ net63 net917 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12735__A cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__C1 _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ net2785 _01996_ net38 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a21o_1
XANTENNA__07388__X _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07997__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13290_ clknet_leaf_23_clk cpu.RU0.next_FetchedInstr\[29\] net1178 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12880__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12241_ cpu.LCD0.row_1\[61\] _06025_ _06027_ cpu.LCD0.row_2\[45\] _06136_ vssd1 vssd1
+ vccd1 vccd1 _06137_ sky130_fd_sc_hd__a221o_1
XANTENNA__09738__A3 _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10202__B1 cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ cpu.LCD0.row_1\[66\] _06001_ _06025_ cpu.LCD0.row_1\[58\] vssd1 vssd1 vccd1
+ vccd1 _06071_ sky130_fd_sc_hd__a22o_1
XANTENNA__07267__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__B1 _02210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net2503 net183 net420 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12470__A cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ net2843 net185 net428 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ cpu.IM0.address_IM\[14\] _05271_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07851__X _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13386__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14631__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_101_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ net2213 net155 net318 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__mux2_1
XANTENNA__07134__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ net723 _05378_ _05823_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a22o_1
X_14675_ net1397 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
X_11887_ net2877 net152 net326 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ cpu.DM0.readdata\[3\] _05030_ net739 vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__mux2_1
X_13626_ clknet_leaf_93_clk _00739_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10769_ net989 net240 vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2_1
X_13557_ clknet_leaf_73_clk _00670_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10864__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12508_ cpu.f0.i\[7\] _05544_ net257 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _06288_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06643__A a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13488_ clknet_leaf_74_clk _00601_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14011__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12439_ net1991 net731 net500 _06243_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12194__B1 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13249__Q a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__A1 _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11695__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ clknet_leaf_88_clk _01222_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14161__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ net448 _03269_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06931_ net954 cpu.RF0.registers\[12\]\[26\] net765 vssd1 vssd1 vccd1 vccd1 _02222_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13729__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14615__RESET_B net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _03044_ net444 _04925_ net443 _03080_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__o32a_1
XFILLER_0_78_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06862_ net1073 net1068 net1066 net1071 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_2_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08601_ cpu.RF0.registers\[4\]\[4\] net678 _03880_ _03881_ _03883_ vssd1 vssd1 vccd1
+ vccd1 _03892_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09581_ _04670_ _04782_ net472 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__mux2_1
X_06793_ _02082_ _02083_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08532_ cpu.RF0.registers\[8\]\[6\] net707 net667 _03809_ _03812_ vssd1 vssd1 vccd1
+ vccd1 _03823_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13879__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12539__B cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload92_A clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ cpu.RF0.registers\[19\]\[8\] net640 _03752_ _03753_ net667 vssd1 vssd1 vccd1
+ vccd1 _03754_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout153_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07414_ net972 cpu.RF0.registers\[14\]\[0\] net763 vssd1 vssd1 vccd1 vccd1 _02705_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13109__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ _03682_ _03683_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ cpu.RF0.registers\[24\]\[3\] net608 _02622_ _02624_ _02628_ vssd1 vssd1 vccd1
+ vccd1 _02636_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__A1 cpu.DM0.readdata\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07276_ net980 cpu.RF0.registers\[6\]\[7\] net802 vssd1 vssd1 vccd1 vccd1 _02567_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10983__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ net1074 cpu.RF0.registers\[29\]\[31\] net848 vssd1 vssd1 vccd1 vccd1 _04306_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13259__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14504__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1327_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 cpu.DM0.readdata\[0\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09864__A cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 cpu.f0.data_adr\[15\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__A1 cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 cpu.RF0.registers\[31\]\[22\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 cpu.RF0.registers\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 cpu.LCD0.row_1\[127\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 cpu.RF0.registers\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 a1.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _02139_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_2
Xfanout621 net624 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_8
Xfanout632 _02100_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlymetal6s2s_1
X_09917_ cpu.IG0.Instr\[27\] net520 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1
+ _05203_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout643 net645 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_8
Xfanout654 net656 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout954_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14654__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout665 _02050_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10499__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 _02039_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09848_ net278 _04442_ _05135_ _05138_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a211o_1
Xfanout687 _02030_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_6
Xfanout698 _02023_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ _05047_ _05048_ _02759_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07390__Y _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ net1816 net210 net335 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__mux2_1
X_12790_ cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08646__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net1549 net219 net342 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__mux2_1
XANTENNA__07550__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14460_ clknet_leaf_23_clk _01570_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11672_ net2328 net229 net352 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ cpu.LCD0.row_1\[29\] cpu.LCD0.row_1\[37\] net896 vssd1 vssd1 vccd1 vccd1
+ _00253_ sky130_fd_sc_hd__mux2_1
X_13411_ clknet_leaf_79_clk _00524_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ clknet_leaf_18_clk _01502_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07559__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ clknet_leaf_42_clk _00455_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_10554_ net1132 net2135 net912 _05664_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__a31o_1
XANTENNA__06463__A a1.WRITE_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12184__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08381__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ clknet_leaf_24_clk cpu.RU0.next_FetchedInstr\[12\] net1205 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[12\] sky130_fd_sc_hd__dfrtp_1
X_10485_ net1448 net922 net747 a1.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__a22o_1
XANTENNA__14184__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12224_ cpu.LCD0.row_2\[92\] _05983_ _06000_ cpu.LCD0.row_2\[60\] vssd1 vssd1 vccd1
+ vccd1 _06121_ sky130_fd_sc_hd__a22o_1
XANTENNA__09774__A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06750__X _02041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10726__A1 a1.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12155_ cpu.LCD0.row_1\[57\] _06025_ _06027_ cpu.LCD0.row_2\[41\] _06054_ vssd1 vssd1
+ vccd1 vccd1 _06055_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11106_ net2697 net248 net421 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__mux2_1
XANTENNA__12479__A1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12086_ cpu.LCD0.nextState\[1\] cpu.LCD0.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05987_
+ sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_88_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__14097__RESET_B net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ net2171 net255 net429 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
XANTENNA__07577__A_N _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07107__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ clknet_leaf_36_clk net1439 net1263 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08556__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11939_ net1939 net218 net318 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14658_ net72 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ clknet_leaf_105_clk _00722_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08607__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14589_ clknet_leaf_49_clk _01691_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[100\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13401__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07130_ _02418_ _02419_ _02420_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10965__A1 _02901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07061_ net1052 cpu.RF0.registers\[17\]\[18\] net806 vssd1 vssd1 vccd1 vccd1 _02352_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12167__B1 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09684__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09032__B1 _04321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13551__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10717__B2 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08240__D1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07963_ cpu.RF0.registers\[12\]\[29\] net697 net685 cpu.RF0.registers\[24\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07635__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_79_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08138__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06914_ cpu.RF0.registers\[8\]\[27\] net611 _02170_ _02174_ _02192_ vssd1 vssd1 vccd1
+ vccd1 _02205_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ _03195_ net448 _04541_ _04986_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a2bb2o_1
X_07894_ cpu.RF0.registers\[22\]\[29\] _02146_ net595 cpu.RF0.registers\[7\]\[29\]
+ _03174_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__a221o_1
XANTENNA__10910__X _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06845_ net1038 cpu.RF0.registers\[23\]\[27\] net817 vssd1 vssd1 vccd1 vccd1 _02136_
+ sky130_fd_sc_hd__and3_1
X_09633_ _03079_ net443 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_84_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09850__C _05131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07651__B _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _04457_ _04460_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06776_ cpu.RF0.registers\[4\]\[30\] net677 net650 cpu.RF0.registers\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14057__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ net1105 cpu.RF0.registers\[29\]\[6\] net849 vssd1 vssd1 vccd1 vccd1 _03806_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08466__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07649__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09495_ _02473_ _03664_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nand2_1
XANTENNA__07370__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ cpu.RF0.registers\[8\]\[8\] net707 net639 cpu.RF0.registers\[26\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ _03664_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07328_ net982 cpu.RF0.registers\[10\]\[3\] net788 vssd1 vssd1 vccd1 vccd1 _02619_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13331__RESET_B net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10517__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__A1 _02543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ net1062 cpu.RF0.registers\[26\]\[7\] net788 vssd1 vssd1 vccd1 vccd1 _02550_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1232_X net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__B1 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ cpu.f0.i\[14\] _05509_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nor2_1
XANTENNA__09023__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__B _03115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _04123_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14190__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
Xfanout473 net477 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
X_13960_ clknet_leaf_99_clk _01073_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout484 _02642_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
Xfanout495 _02089_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
X_12911_ clknet_leaf_25_clk _00100_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13891_ clknet_leaf_78_clk _01004_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12842_ clknet_leaf_31_clk _00061_ net1207 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09105__Y _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12773_ net1460 net496 net281 cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
XANTENNA__13352__Q cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ clknet_leaf_47_clk _01614_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11724_ net1982 net161 net348 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06745__X _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14443_ clknet_leaf_27_clk _01553_ net1188 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_11655_ net1684 net163 net354 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11303__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10606_ cpu.LCD0.row_1\[12\] cpu.LCD0.row_1\[20\] net901 vssd1 vssd1 vccd1 vccd1
+ _00236_ sky130_fd_sc_hd__mux2_1
X_14374_ clknet_leaf_32_clk _01485_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11586_ net1866 net171 net363 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13574__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10537_ net44 net919 vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__and2_1
X_13325_ clknet_leaf_30_clk cpu.RU0.next_dhit net1208 vssd1 vssd1 vccd1 vccd1 cpu.DM0.dhit
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_90_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_4
X_13256_ clknet_leaf_36_clk _00436_ net1264 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10468_ net18 net754 net564 a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06921__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ net743 _05996_ net557 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__and3_1
X_13187_ clknet_leaf_34_clk _00367_ net1245 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10443__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ _01802_ net271 _05617_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06640__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14207__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ _06020_ _06026_ _06032_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11973__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__B cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ cpu.LCD0.cnt_500hz\[11\] _01957_ _05969_ vssd1 vssd1 vccd1 vccd1 _05974_
+ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_1_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09868__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__A1 cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ _01757_ _01968_ _01976_ _01985_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__and4_1
XANTENNA__07471__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06368__A cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__inv_2
XANTENNA__07190__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ cpu.RF0.registers\[28\]\[13\] net705 net684 cpu.RF0.registers\[24\]\[13\]
+ _03569_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09679__A _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09280_ _04569_ _04570_ net455 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__mux2_1
X_06492_ cpu.FetchedInstr\[3\] cpu.FetchedInstr\[2\] _01881_ _01882_ vssd1 vssd1 vccd1
+ vccd1 _01883_ sky130_fd_sc_hd__or4_2
XANTENNA__08583__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08231_ cpu.RF0.registers\[28\]\[14\] net706 net671 cpu.RF0.registers\[23\]\[14\]
+ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a221o_1
XANTENNA__13917__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11213__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ net1099 cpu.RF0.registers\[26\]\[20\] net861 vssd1 vssd1 vccd1 vccd1 _03453_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07199__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07113_ cpu.RF0.registers\[19\]\[14\] net615 net609 cpu.RF0.registers\[3\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ cpu.RF0.registers\[12\]\[22\] net696 net677 cpu.RF0.registers\[4\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22o_1
XANTENNA__12941__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload50 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07044_ cpu.RF0.registers\[8\]\[19\] net611 net584 cpu.RF0.registers\[2\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a22o_1
Xclkload61 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload61/X sky130_fd_sc_hd__clkbuf_4
Xclkload72 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload72/X sky130_fd_sc_hd__clkbuf_4
Xclkload83 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_4
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload94 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__08359__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06550__B net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__C net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _04246_ _04280_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout485_A _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__B2 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net495 _03235_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__xor2_1
X_07877_ _03161_ _03163_ _03165_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10800__B _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13447__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09616_ net458 _04906_ _04905_ _02758_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__o211a_1
X_06828_ _02112_ _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__nor2_1
XANTENNA__08196__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ _02545_ net435 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06759_ net941 net841 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__and2_4
XANTENNA__12567__X _06332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net289 _04765_ _04768_ net297 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08924__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08429_ cpu.RF0.registers\[3\]\[9\] net642 _03702_ _03711_ _03712_ vssd1 vssd1 vccd1
+ vccd1 _03720_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11123__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
X_11440_ net2137 net233 net380 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
XANTENNA__09101__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__A2 _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ net2157 net250 net387 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__mux2_1
XANTENNA__12743__A _06342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ clknet_leaf_54_clk net1806 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_10322_ cpu.f0.i\[21\] net1019 _05549_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14090_ clknet_leaf_101_clk _01203_ net1213 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ clknet_leaf_45_clk _00221_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[5\]
+ sky130_fd_sc_hd__dfstp_1
X_10253_ net1416 _05502_ net725 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14300__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
X_10184_ cpu.IM0.address_IM\[29\] _03193_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nor2_1
XANTENNA__14222__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1213 net1220 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13347__Q cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1224 net1227 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11793__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1235 net1268 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 net1255 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08770__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1257 net1267 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_4
Xfanout1268 net1386 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_4
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout281 _01767_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
Xfanout1279 net1283 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_4
Xfanout292 _04400_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ clknet_leaf_65_clk _01056_ net1282 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14372__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874_ clknet_leaf_70_clk _00987_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12814__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12606__A1 cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ clknet_leaf_14_clk _00044_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12756_ net1586 net497 net279 cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11707_ net2153 net222 net348 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
X_12687_ net2208 cpu.LCD0.row_2\[81\] net1009 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12964__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06635__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14426_ clknet_leaf_17_clk _01537_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11638_ net1912 net234 net356 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11968__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ clknet_leaf_72_clk _01470_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11569_ net2820 net251 net365 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06922__Y _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold707 cpu.RF0.registers\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold718 cpu.RF0.registers\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_16_clk cpu.RU0.next_FetchedData\[15\] net1196 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[15\] sky130_fd_sc_hd__dfrtp_1
Xhold729 a1.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ clknet_leaf_75_clk _01401_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06651__A a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14641__Q cpu.f0.write_data\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ clknet_leaf_37_clk _00419_ net1258 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07185__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07800_ net959 cpu.RF0.registers\[2\]\[22\] net769 vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__and3_1
Xhold1407 a1.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
X_08780_ cpu.RF0.registers\[1\]\[18\] net713 net635 cpu.RF0.registers\[16\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a22o_1
Xhold1418 a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 cpu.K0.code\[4\] vssd1 vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08578__A _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07731_ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__inv_2
XANTENNA__10305__C1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11208__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07662_ net1024 cpu.RF0.registers\[20\]\[16\] net780 vssd1 vssd1 vccd1 vccd1 _02953_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08865__X _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09401_ net449 _04502_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__nand2_1
X_06613_ _01980_ _01981_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__or2_1
X_07593_ net1047 cpu.RF0.registers\[25\]\[12\] net757 vssd1 vssd1 vccd1 vccd1 _02884_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ net474 _04604_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nor2_1
X_06544_ cpu.f0.num\[12\] _01805_ cpu.f0.num\[15\] _01808_ _01914_ vssd1 vssd1 vccd1
+ vccd1 _01933_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ _04205_ _04553_ _03407_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a21oi_1
X_06475_ cpu.K0.code\[4\] cpu.K0.code\[5\] cpu.K0.code\[6\] cpu.K0.code\[7\] vssd1
+ vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__or4b_2
XFILLER_0_5_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10348__A cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08214_ cpu.IM0.address_IM\[21\] net552 _03503_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_
+ sky130_fd_sc_hd__a22o_2
X_09194_ _04483_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__and2_1
XANTENNA__09226__B1 _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10067__B cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11878__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _03434_ _03435_ cpu.IM0.address_IM\[23\] net551 vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA_fanout400_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A0 _03077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07657__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ cpu.RF0.registers\[12\]\[25\] net696 net684 cpu.RF0.registers\[24\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a22o_1
XANTENNA__07252__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14245__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__A1 _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07027_ net1040 cpu.RF0.registers\[21\]\[19\] net796 vssd1 vssd1 vccd1 vccd1 _02318_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10083__A cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__A cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13167__Q a1.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 cpu.RF0.registers\[0\]\[18\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 cpu.f0.write_data\[16\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14395__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 cpu.c0.count\[8\] vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ cpu.RF0.registers\[13\]\[26\] net659 net642 cpu.RF0.registers\[3\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a22o_1
XANTENNA__08488__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold45 _00182_ vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 cpu.f0.data_adr\[20\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 net100 vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 _00164_ vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07929_ cpu.RF0.registers\[18\]\[30\] net580 _03202_ _03207_ _03212_ vssd1 vssd1
+ vccd1 vccd1 _03220_ sky130_fd_sc_hd__a2111o_1
Xhold89 _00162_ vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ net2693 net927 _05676_ net274 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ net723 _05263_ _05797_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12987__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12610_ cpu.LCD0.row_2\[12\] cpu.LCD0.row_2\[4\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13590_ clknet_leaf_58_clk _00703_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06736__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09112__A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__C _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12541_ cpu.K0.code\[4\] cpu.K0.code\[5\] cpu.K0.code\[7\] cpu.K0.code\[6\] vssd1
+ vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or4b_2
XFILLER_0_13_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ net257 _06265_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nor2_1
XANTENNA__07491__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ clknet_leaf_77_clk _01324_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11788__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11024__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ net1809 net167 net383 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XANTENNA__12473__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ clknet_leaf_84_clk _01255_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11354_ net2413 net186 net391 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
XANTENNA__07243__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ net540 _05544_ _05545_ net526 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a211o_1
X_11285_ net1786 net173 net400 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__mux2_1
X_14073_ clknet_leaf_13_clk _01186_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13612__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ clknet_leaf_35_clk _00213_ net1261 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
X_10236_ _01799_ _05482_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_2
Xfanout1021 cpu.f0.i\[7\] vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_4
XANTENNA__09940__A1 cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlymetal6s2s_1
X_10167_ _02004_ _05146_ _05431_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__o211a_1
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_2
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10550__A2 a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1065 net1066 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_2
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_2
X_10098_ cpu.IM0.address_IM\[22\] _03116_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__and2_1
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_1
XANTENNA__09689__A_N _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11028__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ clknet_leaf_5_clk _01039_ net1148 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13857_ clknet_leaf_63_clk _00970_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12808_ clknet_leaf_37_clk _00027_ net1266 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06646__A a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ clknet_leaf_12_clk _00901_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__A1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _01872_ _01763_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09208__A0 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13142__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14268__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14293__RESET_B net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ clknet_leaf_35_clk _01520_ net1258 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09676__B _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07477__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold504 cpu.RF0.registers\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold515 cpu.RF0.registers\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06381__A cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 cpu.RF0.registers\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 cpu.RF0.registers\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold548 cpu.FetchedInstr\[2\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09950_ cpu.IM0.address_IM\[10\] _02474_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__nor2_1
Xhold559 cpu.RF0.registers\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13292__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ _04181_ _04183_ _04188_ _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or4_2
X_09881_ cpu.IM0.address_IM\[3\] net933 _05169_ _05170_ vssd1 vssd1 vccd1 vccd1 _00026_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload18_A clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ _04121_ _04122_ cpu.IM0.address_IM\[19\] net551 vssd1 vssd1 vccd1 vccd1 _04123_
+ sky130_fd_sc_hd__a2bb2o_2
Xhold1204 cpu.RF0.registers\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A0 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 cpu.RF0.registers\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1226 cpu.RF0.registers\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 cpu.RF0.registers\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ _03540_ _03568_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nand3_1
Xhold1248 cpu.LCD0.row_1\[30\] vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 cpu.RF0.registers\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10829__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ net952 cpu.RF0.registers\[2\]\[17\] net769 vssd1 vssd1 vccd1 vccd1 _03005_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ cpu.RF0.registers\[10\]\[1\] net693 net641 cpu.RF0.registers\[19\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_69_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ cpu.RF0.registers\[27\]\[13\] net591 _02916_ _02926_ _02927_ vssd1 vssd1
+ vccd1 vccd1 _02936_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12558__A _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout350_A _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09447__A0 _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _02544_ _02865_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ net485 _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__nor2_1
X_06527_ cpu.f0.num\[4\] _01794_ cpu.f0.num\[14\] _01806_ vssd1 vssd1 vccd1 vccd1
+ _01916_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _04532_ _04536_ net484 vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06458_ _01842_ _01858_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[14\] sky130_fd_sc_hd__and2b_1
XANTENNA__08771__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09177_ net463 _03833_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__nor2_1
X_06389_ cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_78_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13635__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ net1078 cpu.RF0.registers\[21\]\[23\] net866 vssd1 vssd1 vccd1 vccd1 _03419_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08973__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ net943 cpu.RF0.registers\[1\]\[25\] net883 vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__and3_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__06984__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11070_ net1817 net238 net424 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__13785__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ cpu.IM0.address_IM\[16\] _02947_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__nand2_1
XANTENNA__09922__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__C net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12285__A2 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net2188 net218 net314 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
XANTENNA__12739__Y _01767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_83_clk _00824_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10923_ cpu.DM0.readdata\[27\] net734 net719 vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13642_ clknet_leaf_101_clk _00755_ net1213 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10854_ net1588 net224 net432 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
XANTENNA__13165__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10048__A1 cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__Q cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08384__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14410__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ clknet_leaf_9_clk _00686_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ net1823 net559 net538 _05736_ vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08110__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12524_ cpu.f0.i\[26\] _06296_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ cpu.f0.i\[1\] _06250_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06472__Y cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14560__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11406_ net2114 net243 net384 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
X_12386_ net1121 net1533 net530 cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1 vccd1 _01512_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10220__A1 cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10220__B2 cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14125_ clknet_leaf_102_clk _01238_ net1215 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11337_ net1953 net253 net392 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06975__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ clknet_leaf_99_clk _01169_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11268_ cpu.IG0.Instr\[9\] cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__and2b_2
X_13007_ clknet_leaf_35_clk _00196_ net1259 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09913__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ cpu.f0.data_adr\[3\] net729 _05478_ cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1
+ _00056_ sky130_fd_sc_hd__a22o_1
X_11199_ net2754 net143 net412 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__C _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11981__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10287__A1 _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13508__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ clknet_leaf_73_clk _01022_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_07430_ net1056 cpu.RF0.registers\[23\]\[1\] net819 vssd1 vssd1 vccd1 vccd1 _02721_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06376__A cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14090__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07361_ net977 cpu.RF0.registers\[9\]\[2\] net760 vssd1 vssd1 vccd1 vccd1 _02652_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08637__D1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13658__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08101__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ net514 _02112_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__nand2_4
XFILLER_0_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07292_ cpu.IG0.Instr\[11\] net742 _02208_ net1047 vssd1 vssd1 vccd1 vccd1 _02583_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07455__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08591__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ cpu.RF0.registers\[0\]\[31\] net661 net547 vssd1 vssd1 vccd1 vccd1 _04322_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12736__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09601__A0 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07207__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__A2 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 cpu.RF0.registers\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold312 cpu.RF0.registers\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 a1.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold334 cpu.DM0.readdata\[23\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__Y _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__B2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 cpu.RF0.registers\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__X _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold356 cpu.RF0.registers\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold367 cpu.RF0.registers\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold378 cpu.RF0.registers\[16\]\[22\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net717 net134 _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a211oi_1
Xhold389 cpu.RF0.registers\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 _02145_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_4
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_4
Xfanout825 net827 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09904__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08707__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 _02062_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_6
X_09864_ cpu.IM0.address_IM\[0\] _02682_ _05153_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_
+ sky130_fd_sc_hd__and4_1
Xfanout847 _02044_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_6
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_2
XANTENNA__10514__A2 a1.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 cpu.LCD0.row_1\[51\] vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _02016_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 cpu.RF0.registers\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08815_ net938 cpu.RF0.registers\[12\]\[19\] net867 vssd1 vssd1 vccd1 vccd1 _04106_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08469__C net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 cpu.LCD0.row_1\[110\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07373__C net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ _05077_ _05078_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__o21ai_4
Xhold1034 _01710_ vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__A1 cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_A _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 cpu.RF0.registers\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 _00234_ vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__B2 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1067 cpu.LCD0.row_2\[106\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _03836_ _03870_ _04035_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand4_1
XANTENNA__09668__B1 _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__A2 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1078 _01673_ vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06838__X _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 cpu.RF0.registers\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ net1103 cpu.RF0.registers\[27\]\[1\] net881 vssd1 vssd1 vccd1 vccd1 _03968_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1095_X net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ net1036 cpu.RF0.registers\[16\]\[13\] net831 vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13180__Q a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ net1052 cpu.RF0.registers\[30\]\[8\] net763 vssd1 vssd1 vccd1 vccd1 _02850_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1262_X net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10570_ net1132 net1612 net912 _05672_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__a31o_1
XANTENNA__09597__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12735__B _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08932__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ net495 net448 net465 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06733__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12240_ cpu.LCD0.row_1\[45\] _06030_ _06033_ cpu.LCD0.row_2\[77\] vssd1 vssd1 vccd1
+ vccd1 _06136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07548__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A1 cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ cpu.LCD0.row_1\[50\] _06019_ _06037_ cpu.LCD0.row_1\[74\] _06069_ vssd1 vssd1
+ vccd1 vccd1 _06070_ sky130_fd_sc_hd__a221o_1
XANTENNA__08946__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10823__X _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__A1 cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ net1946 net172 net419 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold890 _00235_ vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12470__B cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08159__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ net1926 net190 net426 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XANTENNA__10271__A cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__Y _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10505__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ net715 net133 _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08379__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12258__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07580__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11955_ net2450 net162 net321 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08331__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10906_ cpu.DM0.readdata\[22\] net735 net720 vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__o21a_1
X_14674_ net1396 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__13800__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11886_ net2418 net164 net326 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13625_ clknet_leaf_14_clk _00738_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10837_ net1933 net249 net431 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ clknet_leaf_70_clk _00669_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10768_ a1.ADR_I\[15\] net558 net536 _05724_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__a22o_1
XANTENNA__06924__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08842__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ net1020 _06286_ _06287_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ clknet_leaf_83_clk _00600_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ net2900 cpu.LCD0.row_1\[113\] net906 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XANTENNA__06643__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12438_ cpu.DM0.data_i\[27\] net534 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08398__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11976__S net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12369_ net1121 net1859 net531 cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 _01495_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14306__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14108_ clknet_leaf_11_clk _01221_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06930_ net1029 cpu.RF0.registers\[31\]\[26\] net825 vssd1 vssd1 vccd1 vccd1 _02221_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14039_ clknet_leaf_65_clk _01152_ net1278 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13330__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ net1038 cpu.RF0.registers\[29\]\[27\] net792 vssd1 vssd1 vccd1 vccd1 _02152_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07193__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08600_ cpu.RF0.registers\[11\]\[4\] net688 net657 cpu.RF0.registers\[13\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a22o_1
XANTENNA__08570__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12249__A2 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ net291 _04867_ _04870_ net299 _04869_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a221o_1
X_06792_ cpu.CU0.opcode\[6\] cpu.CU0.opcode\[4\] vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__and2b_2
XANTENNA__08586__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ cpu.RF0.registers\[15\]\[6\] net683 net675 cpu.RF0.registers\[6\]\[6\] _03807_
+ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07921__C net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06377__Y _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13480__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11216__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12539__C cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08462_ net1095 cpu.RF0.registers\[23\]\[8\] net845 vssd1 vssd1 vccd1 vccd1 _03753_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload85_A clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07413_ net1049 cpu.RF0.registers\[30\]\[0\] net763 vssd1 vssd1 vccd1 vccd1 _02704_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08393_ cpu.RF0.registers\[12\]\[10\] net696 net671 cpu.RF0.registers\[23\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout146_A _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ cpu.RF0.registers\[12\]\[3\] net571 _02616_ _02618_ _02629_ vssd1 vssd1 vccd1
+ vccd1 _02635_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_77_clk_X clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07275_ net980 cpu.RF0.registers\[4\]\[7\] net782 vssd1 vssd1 vccd1 vccd1 _02566_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10356__A cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_A _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09014_ net1075 cpu.RF0.registers\[30\]\[31\] net837 vssd1 vssd1 vccd1 vccd1 _04305_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_76_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07368__C net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold120 cpu.FetchedInstr\[3\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09864__B _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 cpu.f0.data_adr\[30\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 cpu.DM0.readdata\[16\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 cpu.RF0.registers\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 cpu.RF0.registers\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _00343_ vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 cpu.RF0.registers\[17\]\[17\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 cpu.RF0.registers\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _02154_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
Xfanout611 _02138_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_6
X_09916_ _05201_ _05202_ cpu.IM0.address_IM\[6\] net933 vssd1 vssd1 vccd1 vccd1 _00029_
+ sky130_fd_sc_hd__a2bb2o_1
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout633 _02084_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
XANTENNA_hold1428_A cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout666 _02050_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_2
X_09847_ _05136_ _05137_ _02437_ net300 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__o2bb2a_1
Xfanout677 _02037_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_6
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 _02028_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_8
Xfanout699 net701 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06568__X _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _04406_ _04966_ _04967_ net299 _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a221o_1
XANTENNA__13823__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08927__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ cpu.RF0.registers\[30\]\[0\] net1096 net839 vssd1 vssd1 vccd1 vccd1 _04020_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11126__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11740_ net2281 net220 net343 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13973__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ net2347 net232 net352 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ clknet_leaf_95_clk _00523_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622_ cpu.LCD0.row_1\[28\] cpu.LCD0.row_1\[36\] net903 vssd1 vssd1 vccd1 vccd1
+ _00252_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07419__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14390_ clknet_leaf_19_clk net1456 net1180 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12412__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__A _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ clknet_leaf_64_clk _00454_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10553_ net53 net919 vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13272_ clknet_leaf_23_clk cpu.RU0.next_FetchedInstr\[11\] net1194 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[11\] sky130_fd_sc_hd__dfrtp_1
X_10484_ net1473 net922 net747 a1.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11796__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ cpu.LCD0.row_2\[124\] _06022_ _06028_ cpu.LCD0.row_1\[116\] _06119_ vssd1
+ vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07575__A _02865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ cpu.LCD0.row_2\[65\] _05988_ _06019_ cpu.LCD0.row_1\[49\] vssd1 vssd1 vccd1
+ vccd1 _06054_ sky130_fd_sc_hd__a22o_1
XANTENNA__13353__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11105_ cpu.RF0.registers\[3\]\[2\] net252 net421 vssd1 vssd1 vccd1 vccd1 _00538_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12479__A2 cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ _05981_ _05984_ net743 vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__and3_4
X_11036_ net1559 net237 net428 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ clknet_leaf_44_clk net1482 net1305 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06638__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11036__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ net1732 net223 net321 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ clknet_leaf_55_clk _01758_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11869_ net1609 net234 net328 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ clknet_leaf_98_clk _00721_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12403__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588_ clknet_leaf_46_clk net2307 net1356 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14644__Q cpu.f0.write_data\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13539_ clknet_leaf_79_clk _00652_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07060_ net1063 cpu.RF0.registers\[18\]\[18\] net771 vssd1 vssd1 vccd1 vccd1 _02351_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07291__B1 _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07188__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12167__B2 cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__A1 cpu.IM0.address_IM\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A2 _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11914__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07485__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07916__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ cpu.RF0.registers\[22\]\[29\] net670 net649 cpu.RF0.registers\[14\]\[29\]
+ _03245_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a221o_1
XANTENNA__13846__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _04912_ _04360_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand2b_1
X_06913_ cpu.RF0.registers\[10\]\[27\] net569 _02149_ _02136_ net624 vssd1 vssd1 vccd1
+ vccd1 _02204_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ cpu.RF0.registers\[2\]\[29\] net585 _02195_ cpu.RF0.registers\[30\]\[29\]
+ _03183_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09632_ _03079_ net443 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06844_ net1039 net817 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06829__A _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__D _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09205__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12870__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _04770_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__nand2_1
XANTENNA__13996__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06775_ net1089 net841 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_65_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06548__B net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ net949 cpu.RF0.registers\[7\]\[6\] net846 vssd1 vssd1 vccd1 vccd1 _03805_
+ sky130_fd_sc_hd__and3_1
X_09494_ _02473_ _03664_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__or2_1
XANTENNA__07649__A2 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ cpu.RF0.registers\[1\]\[8\] net713 net643 cpu.RF0.registers\[3\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09859__B _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout430_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13226__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ _02473_ _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_22_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08482__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07327_ net975 cpu.RF0.registers\[13\]\[3\] net793 vssd1 vssd1 vccd1 vccd1 _02618_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08074__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07098__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13376__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ net980 cpu.RF0.registers\[1\]\[7\] net806 vssd1 vssd1 vccd1 vccd1 _02549_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07821__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__B2 cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07189_ net1046 cpu.RF0.registers\[23\]\[10\] net817 vssd1 vssd1 vccd1 vccd1 _02480_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 net433 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 _04086_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout452 _02757_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_2
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net477 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout485 _02642_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout496 _01761_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
X_12910_ clknet_leaf_26_clk _00099_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07888__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ clknet_leaf_11_clk _01003_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09115__A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08657__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14001__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ clknet_leaf_30_clk _00060_ net1207 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07561__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ net1467 net496 net281 cpu.f0.i\[30\] vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08954__A _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ clknet_leaf_55_clk net2498 net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11723_ net2065 net178 net347 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14151__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14442_ clknet_leaf_27_clk _01552_ net1183 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_11654_ net2020 net169 net355 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
XANTENNA__06474__A cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12397__A1 cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13719__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14464__Q cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ net2295 cpu.LCD0.row_1\[19\] net899 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06905__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14373_ clknet_leaf_32_clk _01484_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08065__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ net2159 net186 net364 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__mux2_1
Xwire842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ clknet_leaf_17_clk cpu.RU0.next_FetchedData\[31\] net1194 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[31\] sky130_fd_sc_hd__dfrtp_1
X_10536_ net1134 net2872 net914 _05655_ vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_90_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06761__X _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_23_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ clknet_leaf_21_clk _00435_ net1171 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06480__Y _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ net17 net752 net562 net1712 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__o22a_1
XANTENNA__13869__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__B _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ net745 _06009_ _06014_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or4_1
X_13186_ clknet_leaf_34_clk _00366_ net1208 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10443__B net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ net1124 _01803_ net267 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or3_1
X_12137_ cpu.LCD0.row_1\[16\] _06036_ _06037_ cpu.LCD0.row_1\[72\] _06035_ vssd1 vssd1
+ vccd1 vccd1 _06038_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12893__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ _05973_ net502 _05972_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__and3b_1
XANTENNA__14247__RESET_B net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ cpu.f0.write_data\[28\] _05898_ net993 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__mux2_1
XANTENNA__07752__B _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14639__Q cpu.f0.write_data\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13249__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ net988 cpu.f0.write_i _01943_ _01780_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06491_ cpu.FetchedInstr\[0\] cpu.FetchedInstr\[1\] vssd1 vssd1 vccd1 vccd1 _01882_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09679__B _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07500__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ cpu.RF0.registers\[11\]\[14\] net688 net639 cpu.RF0.registers\[26\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13882__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13399__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__A1_N net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12388__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14644__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__B2 cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08161_ _03448_ _03449_ _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07112_ cpu.RF0.registers\[6\]\[14\] net583 net565 cpu.RF0.registers\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09695__A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ net936 cpu.RF0.registers\[14\]\[22\] net837 vssd1 vssd1 vccd1 vccd1 _03383_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_41_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload40 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_6
X_07043_ net1040 cpu.RF0.registers\[28\]\[19\] net766 vssd1 vssd1 vccd1 vccd1 _02334_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkload48_A clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload51 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload62 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__bufinv_16
Xclkload73 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_6
Xclkload84 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__clkinv_4
Xclkload95 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12560__B2 _06326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__inv_2
XANTENNA__09308__A2 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14024__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A _03233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ net495 _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07876_ cpu.RF0.registers\[23\]\[28\] net613 net607 cpu.RF0.registers\[24\]\[28\]
+ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a221o_1
XANTENNA__07724__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ net463 _03964_ _04464_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__o21ba_1
X_06827_ _02115_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout645_A _02063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09546_ _02544_ _03729_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__or2_1
X_06758_ net1114 net1116 net1110 net1112 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__nor4_2
XANTENNA__08774__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09477_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__inv_2
XANTENNA__08295__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout812_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06689_ net1858 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[25\] sky130_fd_sc_hd__and2_1
XANTENNA__11404__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08428_ cpu.RF0.registers\[24\]\[9\] net684 net636 cpu.RF0.registers\[16\]\[9\] _03703_
+ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload1 clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08359_ cpu.RF0.registers\[31\]\[11\] net686 net640 cpu.RF0.registers\[19\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__B1_N net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1342_X net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ net2522 net253 net387 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__mux2_1
X_10321_ cpu.f0.i\[21\] net540 _05549_ net1019 vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ clknet_leaf_45_clk _00220_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ net528 _05500_ _05501_ net308 _05499_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a32o_1
XANTENNA__08014__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ cpu.IM0.address_IM\[28\] net932 _05446_ _05447_ vssd1 vssd1 vccd1 vccd1 _00051_
+ sky130_fd_sc_hd__a22o_1
Xfanout1203 net1210 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_2
Xfanout1214 net1220 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
Xfanout1225 net1227 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07853__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1247 net1255 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1258 net1261 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_4
Xfanout260 _06252_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout271 _05604_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06781__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1269 net1272 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__clkbuf_4
Xfanout282 _05868_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
X_13942_ clknet_leaf_59_clk _01055_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14517__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14459__Q cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ clknet_leaf_76_clk _00986_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12824_ clknet_leaf_14_clk _00043_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13541__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ net1441 net496 net281 cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11314__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ net2298 net227 net347 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12686_ net2359 cpu.LCD0.row_2\[80\] net1010 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
X_14425_ clknet_leaf_17_clk _01536_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08038__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11637_ net1847 net242 net356 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
XANTENNA__09011__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14356_ clknet_leaf_72_clk _01469_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06932__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ net2637 net254 net365 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13307_ clknet_leaf_31_clk cpu.RU0.next_FetchedData\[14\] net1205 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08850__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold708 cpu.RF0.registers\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ net66 net918 vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold719 cpu.RF0.registers\[29\]\[28\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ clknet_leaf_82_clk _01400_ net1285 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ cpu.RF0.registers\[14\]\[31\] net128 net374 vssd1 vssd1 vccd1 vccd1 _00919_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06651__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ clknet_leaf_37_clk _00418_ net1264 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14047__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11984__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ clknet_leaf_36_clk _00349_ net1263 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08210__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1408 cpu.K0.code\[1\] vssd1 vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 cpu.RF0.registers\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13071__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _02348_ _02384_ _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or3b_2
XANTENNA__14197__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ net953 cpu.RF0.registers\[9\]\[16\] net756 vssd1 vssd1 vccd1 vccd1 _02952_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ net453 _04506_ _04690_ net301 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06612_ _01980_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ net964 cpu.RF0.registers\[6\]\[12\] _02145_ vssd1 vssd1 vccd1 vccd1 _02883_
+ sky130_fd_sc_hd__and3_1
X_09331_ _02250_ net435 net289 _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o211a_1
X_06543_ cpu.f0.num\[6\] _01797_ _01800_ cpu.f0.i\[10\] _01931_ vssd1 vssd1 vccd1
+ vccd1 _01932_ sky130_fd_sc_hd__a221o_1
XANTENNA__11224__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _04203_ _04210_ _03512_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a21o_1
XANTENNA__11281__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06474_ cpu.DM0.dhit net1128 vssd1 vssd1 vccd1 vccd1 cpu.f0.next_lcd_en sky130_fd_sc_hd__and2_1
XFILLER_0_69_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08213_ cpu.RF0.registers\[0\]\[21\] net662 net548 vssd1 vssd1 vccd1 vccd1 _03504_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ net473 net437 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__nand2_1
XANTENNA__08029__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10916__X _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09777__A2 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ cpu.RF0.registers\[0\]\[23\] net661 net547 vssd1 vssd1 vccd1 vccd1 _03435_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__12230__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__A_N net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ cpu.RF0.registers\[4\]\[25\] _02037_ net642 cpu.RF0.registers\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1135_A _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10792__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07026_ net1040 cpu.RF0.registers\[18\]\[19\] net770 vssd1 vssd1 vccd1 vccd1 _02317_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07376__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__A1 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B _02606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1302_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 cpu.f0.data_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ cpu.RF0.registers\[18\]\[26\] net680 net672 cpu.RF0.registers\[29\]\[26\]
+ _04257_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a221o_1
Xhold24 cpu.f0.write_data\[17\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 cpu.f0.write_data\[13\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 cpu.f0.write_data\[22\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ cpu.RF0.registers\[17\]\[30\] net605 net596 cpu.RF0.registers\[7\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__a22o_1
Xhold57 cpu.RF0.registers\[0\]\[3\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _00157_ vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold79 net86 vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13564__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__Q a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ net488 _02213_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10870_ cpu.DM0.readdata\[12\] net736 net720 vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08935__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ _03471_ _03505_ net441 net440 net461 net454 vssd1 vssd1 vccd1 vccd1 _04820_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08268__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ net1128 cpu.f0.state\[3\] cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 _06308_
+ sky130_fd_sc_hd__or3_2
XANTENNA__09112__B _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ cpu.f0.i\[6\] _06262_ net261 vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__o21ai_1
X_14210_ clknet_leaf_94_clk _01323_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11422_ net2864 net182 net384 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11024__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__B1 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14141_ clknet_leaf_67_clk _01254_ net1294 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11353_ net2387 net189 net390 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14592__RESET_B net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ net1020 _05539_ net308 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__o21ai_1
X_14072_ clknet_leaf_18_clk _01185_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ net2769 net193 net400 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__mux2_1
XANTENNA__13358__Q cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ clknet_leaf_36_clk _00212_ net1264 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13094__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10235_ _01799_ _05482_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__nor2_1
XANTENNA__07854__Y _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 net1012 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_2
XANTENNA__07583__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1022 net1023 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
Xfanout1033 net1037 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
X_10166_ _05428_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a21o_1
XANTENNA__13907__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
Xfanout1055 net1059 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11309__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1066 cpu.IG0.Instr\[23\] vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12288__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1077 net1091 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_2
Xfanout1088 net1090 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_2
X_10097_ _05367_ _05368_ cpu.IM0.address_IM\[21\] net1022 vssd1 vssd1 vccd1 vccd1
+ _00044_ sky130_fd_sc_hd__o2bb2a_1
Xfanout1099 net1108 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XANTENNA__10838__A1 _05030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13925_ clknet_leaf_3_clk _01038_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09006__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08900__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12931__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ clknet_leaf_9_clk _00969_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06927__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ clknet_leaf_38_clk _00026_ net1266 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08259__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13787_ clknet_leaf_13_clk _00900_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10999_ _03115_ net532 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__nor2_1
XANTENNA__06646__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ cpu.f0.write_data\[2\] net498 _01762_ _01766_ vssd1 vssd1 vccd1 vccd1 _01723_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11979__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10883__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09208__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ net2141 cpu.LCD0.row_2\[63\] net1002 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__mux2_1
X_14408_ clknet_leaf_35_clk _01519_ net1258 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11015__A1 _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06662__A a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08580__C _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12763__A1 cpu.f0.write_data\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ clknet_leaf_48_clk _01452_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12763__B2 cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10184__A cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold505 cpu.RF0.registers\[21\]\[30\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10774__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 cpu.RF0.registers\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08431__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 cpu.RF0.registers\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold538 cpu.RF0.registers\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09973__A cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 cpu.RF0.registers\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07196__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08900_ cpu.RF0.registers\[18\]\[17\] net680 net665 _04189_ _04190_ vssd1 vssd1 vccd1
+ vccd1 _04191_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12603__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _02101_ _05030_ net1022 vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__o21a_1
XANTENNA__08589__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__B1 _04682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ cpu.RF0.registers\[0\]\[19\] net662 net547 vssd1 vssd1 vccd1 vccd1 _04122_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__06601__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13587__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1205 cpu.RF0.registers\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 cpu.LCD0.row_2\[30\] vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11219__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__B1 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ _03600_ _03630_ _03631_ _03598_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__o31ai_1
Xhold1227 cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 cpu.LCD0.row_1\[87\] vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _00254_ vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ net956 cpu.RF0.registers\[4\]\[17\] net780 vssd1 vssd1 vccd1 vccd1 _03004_
+ sky130_fd_sc_hd__and3_1
X_08693_ _03978_ _03979_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__or3_1
XANTENNA__08498__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout176_A _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07644_ cpu.RF0.registers\[1\]\[13\] net588 _02912_ _02919_ _02923_ vssd1 vssd1 vccd1
+ vccd1 _02935_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07575_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__inv_2
XANTENNA__09447__A1 _03436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _04603_ _04604_ net473 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__mux2_1
X_06526_ cpu.f0.num\[2\] _01792_ cpu.f0.num\[17\] _01810_ vssd1 vssd1 vccd1 vccd1
+ _01915_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14212__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11889__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ _04533_ _04534_ net476 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__mux2_2
XFILLER_0_8_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06457_ cpu.c0.count\[13\] _01843_ cpu.c0.count\[14\] vssd1 vssd1 vccd1 vccd1 _01858_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1252_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__A1 _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07668__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ net468 _03866_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06388_ cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12754__A1 cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__X _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ net1078 cpu.RF0.registers\[29\]\[23\] net848 vssd1 vssd1 vccd1 vccd1 _03418_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_47_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14362__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09883__A cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ net943 cpu.RF0.registers\[8\]\[25\] net873 vssd1 vssd1 vccd1 vccd1 _03349_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__A2 _02271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
X_07009_ cpu.RF0.registers\[9\]\[23\] net573 _02276_ _02278_ _02285_ vssd1 vssd1 vccd1
+ vccd1 _02300_ sky130_fd_sc_hd__a2111o_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
X_10020_ _05296_ _05297_ cpu.IM0.address_IM\[15\] net930 vssd1 vssd1 vccd1 vccd1 _00038_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09922__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__Q cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11129__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07690__X _02981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ net1932 net220 net316 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ clknet_leaf_2_clk _00823_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10922_ net738 _04601_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ clknet_leaf_105_clk _00754_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10853_ net723 _05211_ _05784_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__a22o_4
XANTENNA__09438__A1 _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ clknet_leaf_96_clk _00685_ net1231 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10784_ cpu.IM0.address_IM\[20\] net1014 net285 _05735_ vssd1 vssd1 vccd1 vccd1 _05736_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08962__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11799__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ cpu.f0.i\[25\] _06294_ _06297_ net260 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ _06250_ net263 _06253_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__and3b_1
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14472__Q cpu.SR1.char_in\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11405_ net2819 net245 net384 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12385_ net1119 net1885 net529 cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 _01511_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10756__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14124_ clknet_leaf_87_clk _01237_ net1287 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11336_ net1923 net238 net392 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ clknet_leaf_82_clk _01168_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11267_ net2282 net130 net402 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__mux2_1
XANTENNA__10508__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006_ clknet_leaf_43_clk _00195_ net1303 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
X_10218_ cpu.f0.data_adr\[2\] net729 _05478_ cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _00055_ sky130_fd_sc_hd__a22o_1
XANTENNA__09913__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ net2553 net146 net413 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XANTENNA__13816__Q cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11039__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10149_ cpu.IM0.address_IM\[26\] _02248_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_6_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10878__S _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ clknet_leaf_71_clk _01021_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14235__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ clknet_leaf_83_clk _00952_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07360_ net976 cpu.RF0.registers\[10\]\[2\] net788 vssd1 vssd1 vccd1 vccd1 _02651_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_18_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07291_ net545 _02579_ _02580_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14385__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11502__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ net665 _04313_ _04317_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__or4_2
XFILLER_0_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07860__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07919__C net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__A1 _06326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14382__Q cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__B2 cpu.f0.write_data\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold302 cpu.RF0.registers\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold313 cpu.RF0.registers\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 cpu.RF0.registers\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold335 cpu.RF0.registers\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 cpu.c0.count\[4\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload30_A clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold357 cpu.RF0.registers\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _05214_ _05215_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__and2_1
Xhold368 cpu.RF0.registers\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12977__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold379 cpu.RF0.registers\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout826 net827 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09904__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _01786_ _02719_ _02720_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nand3_1
Xfanout837 _02052_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08112__A _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _02029_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_6
Xhold1002 cpu.RF0.registers\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ net1083 cpu.RF0.registers\[30\]\[19\] net837 vssd1 vssd1 vccd1 vccd1 _04105_
+ sky130_fd_sc_hd__and3_1
Xhold1013 cpu.RF0.registers\[1\]\[28\] vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ net278 _04478_ _05081_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a211oi_2
Xhold1024 _00326_ vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 cpu.LCD0.row_1\[47\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07951__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 cpu.LCD0.row_2\[94\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _03833_ _03835_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__or2_1
Xhold1057 cpu.DM0.readdata\[17\] vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A1 _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 cpu.LCD0.row_2\[113\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 cpu.RF0.registers\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08676_ _03966_ _03964_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07143__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08485__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ net1037 cpu.RF0.registers\[31\]\[13\] net827 vssd1 vssd1 vccd1 vccd1 _02918_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__A cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13602__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07558_ net970 cpu.RF0.registers\[15\]\[8\] net830 vssd1 vssd1 vccd1 vccd1 _02849_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06854__X _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06509_ cpu.f0.num\[1\] cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ net1056 cpu.RF0.registers\[27\]\[5\] net778 vssd1 vssd1 vccd1 vccd1 _02780_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1255_X net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11412__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _03302_ _04289_ _04292_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14184__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09159_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12170_ cpu.LCD0.row_1\[10\] _05994_ _06028_ cpu.LCD0.row_1\[114\] vssd1 vssd1 vccd1
+ vccd1 _06069_ sky130_fd_sc_hd__a22o_1
XANTENNA__10202__A2 _05443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ cpu.RF0.registers\[3\]\[18\] net188 net421 vssd1 vssd1 vccd1 vccd1 _00554_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06811__D1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14108__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 cpu.RF0.registers\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold891 cpu.RF0.registers\[5\]\[0\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ net2367 net207 net426 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
XANTENNA__08022__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10271__B cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07906__A1 _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _05278_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_53_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13132__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11954_ net2372 net178 net320 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14467__Q cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ net735 _04617_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nand2_1
X_14673_ net1395 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
X_11885_ net1675 net168 net327 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13282__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13624_ clknet_leaf_7_clk _00737_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ _01785_ _05773_ net721 vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__mux2_8
XFILLER_0_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13555_ clknet_leaf_67_clk _00668_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10767_ net284 _05722_ _05723_ net1013 cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1
+ vccd1 _05724_ sky130_fd_sc_hd__a32o_1
XANTENNA__10286__X _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11322__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ net1020 _06286_ net262 vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07842__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13486_ clknet_leaf_1_clk _00599_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ cpu.LCD0.row_1\[104\] net2759 net909 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12437_ net2542 net730 net500 _06242_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__o22a_1
XANTENNA__12194__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12368_ net1120 net1646 net530 cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 _01494_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06940__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107_ clknet_leaf_92_clk _01220_ net1241 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11319_ net2912 net206 net394 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
XANTENNA__07755__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net1378 _06191_ _06192_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_97_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14038_ clknet_leaf_71_clk _01151_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07474__C net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ net1049 net793 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06791_ cpu.CU0.opcode\[3\] cpu.CU0.opcode\[2\] cpu.CU0.opcode\[1\] cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__and4b_2
XFILLER_0_54_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08530_ _03818_ _03819_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__or3_1
XANTENNA__13625__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08461_ net1095 cpu.RF0.registers\[24\]\[8\] net871 vssd1 vssd1 vccd1 vccd1 _03752_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07412_ cpu.RF0.registers\[25\]\[0\] net568 _02700_ _02701_ _02702_ vssd1 vssd1 vccd1
+ vccd1 _02703_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_63_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08392_ cpu.RF0.registers\[6\]\[10\] net676 _03675_ _03676_ _03679_ vssd1 vssd1 vccd1
+ vccd1 _03683_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_58_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload78_A clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07343_ cpu.RF0.registers\[9\]\[3\] net573 _02609_ _02615_ _02627_ vssd1 vssd1 vccd1
+ vccd1 _02634_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09822__A1 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_A _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07833__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ net981 cpu.RF0.registers\[9\]\[7\] net759 vssd1 vssd1 vccd1 vccd1 _02565_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09013_ net1074 cpu.RF0.registers\[28\]\[31\] net867 vssd1 vssd1 vccd1 vccd1 _04304_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10924__X _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 net84 vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 net97 vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 cpu.SR1.char_in\[5\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06850__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_1_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 cpu.RF0.registers\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 cpu.RF0.registers\[26\]\[11\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 cpu.RF0.registers\[26\]\[10\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 cpu.LCD0.row_1\[120\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 cpu.FetchedInstr\[12\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _02151_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_8
Xhold198 a1.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13155__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout612 _02138_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_8
X_09915_ _02101_ _04896_ cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o21ai_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout634 _02084_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_42_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14400__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _02063_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_4
Xfanout656 _02056_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10499__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _02436_ net435 _04945_ net293 net289 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__o221a_1
Xfanout667 _02050_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_6
Xfanout678 _02037_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08777__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 _02028_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_2
X_09777_ _02794_ _03866_ _04396_ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a31o_1
X_06989_ net955 cpu.RF0.registers\[14\]\[23\] net761 vssd1 vssd1 vccd1 vccd1 _02280_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11407__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08728_ cpu.RF0.registers\[1\]\[0\] net946 net884 vssd1 vssd1 vccd1 vccd1 _04019_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ cpu.RF0.registers\[13\]\[2\] net657 _03947_ _03948_ _03949_ vssd1 vssd1 vccd1
+ vccd1 _03950_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10120__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11670_ net2620 net244 net352 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10621_ net2303 cpu.LCD0.row_1\[35\] net899 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10959__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11142__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ clknet_leaf_15_clk _00453_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10552_ net1133 net1823 net913 _05663_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__a31o_1
XANTENNA__07285__D1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08017__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13271_ clknet_leaf_23_clk cpu.RU0.next_FetchedInstr\[10\] net1178 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[10\] sky130_fd_sc_hd__dfrtp_1
X_10483_ net1523 net922 net747 a1.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12222_ cpu.LCD0.row_2\[116\] _06007_ _06025_ cpu.LCD0.row_1\[60\] vssd1 vssd1 vccd1
+ vccd1 _06119_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06760__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12153_ cpu.LCD0.row_1\[41\] _06030_ _06037_ cpu.LCD0.row_1\[73\] _06052_ vssd1 vssd1
+ vccd1 vccd1 _06053_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11104_ net2579 net254 net421 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__mux2_1
X_12084_ cpu.LCD0.nextState\[5\] cpu.LCD0.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05985_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__14080__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__X _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _05907_ net504 _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__and3_4
XANTENNA__12701__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13648__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__X _02050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__Y _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12986_ clknet_leaf_28_clk net1501 net1190 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08304__A1 _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09014__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ net1957 net224 net320 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11868_ net2083 net243 net328 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__mux2_1
X_14656_ clknet_leaf_55_clk _01757_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06935__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ net2933 net558 net536 _05760_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__a22o_1
X_13607_ clknet_leaf_78_clk _00720_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13028__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587_ clknet_leaf_54_clk net2248 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_11799_ net2823 net253 net337 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__B2 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13538_ clknet_leaf_94_clk _00651_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11987__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07291__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ clknet_leaf_87_clk _00582_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10891__S net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12167__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13178__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__X _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10717__A3 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ net948 cpu.RF0.registers\[7\]\[29\] net845 vssd1 vssd1 vccd1 vccd1 _03252_
+ sky130_fd_sc_hd__and3_1
X_09700_ _04921_ _04944_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__or2_1
X_06912_ _02199_ _02200_ _02201_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__or4_1
XANTENNA__14573__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ cpu.RF0.registers\[20\]\[29\] _02160_ net587 cpu.RF0.registers\[4\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09740__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ _04608_ _04609_ _04558_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__o21ai_1
X_06843_ net1066 net1068 net1070 net1073 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11227__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ net482 _04741_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06774_ net1092 net861 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08513_ net1102 cpu.RF0.registers\[18\]\[6\] net853 vssd1 vssd1 vccd1 vccd1 _03804_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07006__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _04671_ _04783_ net480 vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout256_A _05772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08444_ _03732_ _03734_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14484__D net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _02508_ _02832_ _02867_ net491 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ net1062 cpu.RF0.registers\[27\]\[3\] net778 vssd1 vssd1 vccd1 vccd1 _02617_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11897__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ net982 cpu.RF0.registers\[5\]\[7\] net797 vssd1 vssd1 vccd1 vccd1 _02548_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1332_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09023__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07188_ net968 cpu.RF0.registers\[12\]\[10\] net766 vssd1 vssd1 vccd1 vccd1 _02479_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_42_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10169__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08231__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08642__A1_N net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout420 _05914_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_6
XFILLER_0_79_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 _03594_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 _02718_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_2
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 _02642_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
Xfanout497 net499 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
X_09829_ _04756_ _04773_ _04846_ _05075_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__or4_1
XANTENNA__13940__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_30_clk _00059_ net1208 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09115__B _04405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ cpu.f0.write_data\[29\] net498 net279 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1
+ _01750_ sky130_fd_sc_hd__a22o_1
XANTENNA__08298__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ clknet_leaf_45_clk _01612_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[21\]
+ sky130_fd_sc_hd__dfstp_1
X_11722_ net2751 net152 net346 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06755__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ clknet_leaf_27_clk _01551_ net1183 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_11653_ net2804 net182 net356 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ net2461 cpu.LCD0.row_1\[18\] net898 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ clknet_leaf_26_clk _01483_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.K0.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ net1592 net191 net362 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14446__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire843 _02049_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
X_13323_ clknet_leaf_16_clk cpu.RU0.next_FetchedData\[30\] net1195 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[30\] sky130_fd_sc_hd__dfrtp_1
X_10535_ net43 net918 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11600__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07586__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire887 _02006_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_2
X_13254_ clknet_leaf_22_clk _00434_ net1171 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net16 net752 net562 net2073 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12205_ _06011_ _06016_ _06021_ _06025_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ clknet_leaf_35_clk _00365_ net1259 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_61_clk_X clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14596__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _01800_ net270 _05616_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13470__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ _05984_ net743 _05989_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and3_4
XFILLER_0_27_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09009__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__A1 cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ cpu.LCD0.cnt_500hz\[9\] cpu.LCD0.cnt_500hz\[10\] _05969_ vssd1 vssd1 vccd1
+ vccd1 _05973_ sky130_fd_sc_hd__and3_1
X_11018_ _03169_ _05847_ net283 vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08848__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08289__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ clknet_leaf_44_clk net1449 net1303 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08828__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10096__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06490_ cpu.FetchedInstr\[4\] cpu.FetchedInstr\[7\] cpu.FetchedInstr\[6\] cpu.FetchedInstr\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_16_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06665__A a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08583__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639_ clknet_leaf_24_clk _01740_ net1210 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09789__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ cpu.RF0.registers\[31\]\[20\] net686 net655 cpu.RF0.registers\[2\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a22o_1
XANTENNA__07249__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_X clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07199__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07111_ _02398_ _02399_ _02400_ _02401_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ net1081 cpu.RF0.registers\[31\]\[22\] net859 vssd1 vssd1 vccd1 vccd1 _03382_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09695__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10915__A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09187__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__13813__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload41 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_6
X_07042_ net962 cpu.RF0.registers\[11\]\[19\] net779 vssd1 vssd1 vccd1 vccd1 _02333_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload52 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload52/X sky130_fd_sc_hd__clkbuf_4
Xclkload63 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_clkbuf_leaf_29_clk_X clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload74 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14390__Q cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload85 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08213__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload96 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__10020__B1 cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _04278_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__and2_2
XANTENNA__13963__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _03198_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07662__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ cpu.RF0.registers\[21\]\[28\] net593 net571 cpu.RF0.registers\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a22o_1
X_09614_ _04472_ _04901_ net458 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o21ai_1
X_06826_ _02102_ _02105_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__o21bai_2
XANTENNA__14319__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _04722_ _04835_ net480 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__mux2_1
X_06757_ net1080 cpu.RF0.registers\[22\]\[30\] net851 vssd1 vssd1 vccd1 vccd1 _02048_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08819__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1282_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _02940_ net442 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06688_ a1.CPU_DAT_O\[24\] net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__14469__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ _03715_ _03716_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ cpu.RF0.registers\[4\]\[11\] net678 _03636_ _03639_ _03642_ vssd1 vssd1 vccd1
+ vccd1 _03649_ sky130_fd_sc_hd__a2111o_1
Xclkload2 clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_8
XANTENNA__12583__Y _06345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07309_ cpu.RF0.registers\[28\]\[4\] net577 _02599_ net622 vssd1 vssd1 vccd1 vccd1
+ _02600_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08289_ cpu.RF0.registers\[18\]\[13\] net680 net659 cpu.RF0.registers\[13\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1335_X net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13493__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10825__A cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11420__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10320_ net2897 _05559_ net724 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__Q cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ cpu.f0.i\[11\] net540 vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__or2_1
XANTENNA__08204__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__A2 cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net630 _04715_ net932 vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a21oi_1
Xfanout1204 net1206 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07022__A4 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1215 net1220 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_2
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_2
Xfanout1237 net1241 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
Xfanout250 _05774_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1248 net1255 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_2
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_2
Xfanout261 _06252_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_1
Xfanout272 _04564_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout283 _05868_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
X_13941_ clknet_leaf_68_clk _01054_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout294 _04397_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13872_ clknet_leaf_76_clk _00985_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08965__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ clknet_leaf_40_clk _00042_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_12754_ cpu.f0.write_data\[12\] net497 net280 cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1
+ _01733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ net1989 net228 net347 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
X_12685_ net2810 net2251 net1002 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XANTENNA__08691__B1 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13836__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ net2093 net245 net356 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
X_14424_ clknet_leaf_17_clk _01535_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06772__X _02063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11567_ net2021 net238 net364 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
X_14355_ clknet_leaf_58_clk _01468_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11330__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ net1135 a1.ADR_I\[3\] net915 _05646_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__a31o_1
X_13306_ clknet_leaf_31_clk cpu.RU0.next_FetchedData\[13\] net1205 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[13\] sky130_fd_sc_hd__dfrtp_1
X_14286_ clknet_leaf_1_clk _01399_ net1142 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 cpu.RF0.registers\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ net2354 net139 net374 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__mux2_1
XANTENNA__12860__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13986__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ clknet_leaf_27_clk _00417_ net1183 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10449_ net29 net755 net564 a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08699__X _03990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ clknet_leaf_36_clk _00348_ net1263 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12119_ cpu.LCD0.row_2\[96\] _06018_ _06019_ cpu.LCD0.row_1\[48\] _06017_ vssd1 vssd1
+ vccd1 vccd1 _06020_ sky130_fd_sc_hd__a221o_1
XANTENNA__13216__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ clknet_leaf_46_clk _00279_ net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1409 cpu.RF0.registers\[16\]\[2\] vssd1 vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07482__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ net1025 cpu.RF0.registers\[17\]\[16\] net804 vssd1 vssd1 vccd1 vccd1 _02951_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07182__B1 _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07721__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ _01757_ _01756_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__xnor2_1
X_07591_ net968 cpu.RF0.registers\[9\]\[12\] net757 vssd1 vssd1 vccd1 vccd1 _02882_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14611__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ net297 net294 _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__mux2_1
X_06542_ _01898_ _01899_ _01908_ _01909_ _01911_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a221o_1
XANTENNA__14385__Q cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _04203_ _04210_ _03477_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06473_ a1.WRITE_I _01789_ a1.curr_state\[0\] net1135 net2414 vssd1 vssd1 vccd1 vccd1
+ _00010_ sky130_fd_sc_hd__a32o_1
XANTENNA__08682__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ _03493_ _03495_ _03500_ _03502_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__or4_1
X_09192_ net449 net437 vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload60_A clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _03430_ net661 _03426_ _03433_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__and4b_1
XFILLER_0_12_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09777__A3 _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_A _05790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ cpu.RF0.registers\[5\]\[25\] net702 net638 cpu.RF0.registers\[26\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a22o_1
XANTENNA__08115__A _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07657__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10792__B2 cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ cpu.RF0.registers\[0\]\[19\] net617 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__or2_1
XANTENNA__09529__A3 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1030_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 net123 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__A cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14141__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _04263_ _04264_ _04265_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__or4_1
Xhold25 cpu.LCD0.row_2\[126\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07018__X _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 cpu.c0.count\[0\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 net95 vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ cpu.RF0.registers\[19\]\[30\] net616 _03211_ _03213_ _03216_ vssd1 vssd1
+ vccd1 vccd1 _03218_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13709__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 cpu.LCD0.row_2\[120\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ net488 _02250_ _03148_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__o21a_1
XANTENNA__06857__X _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ _01999_ _02082_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14291__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06920__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13859__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ _04383_ _04630_ _04815_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_39_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10539__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12808__Q cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _04707_ _04709_ net477 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08673__B1 _03962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__C1 cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10480__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ cpu.f0.i\[5\] cpu.f0.i\[6\] _06260_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12883__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ net1796 net171 net383 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XANTENNA__11150__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10232__B1 _05484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ clknet_leaf_12_clk _01253_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12772__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ net2356 _05810_ net390 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08025__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__A1 _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net540 _05539_ net1020 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13239__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14071_ clknet_leaf_65_clk _01184_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10842__X _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283_ net2757 net197 net398 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__mux2_1
X_13022_ clknet_leaf_34_clk _00211_ net1250 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
X_10234_ cpu.f0.i\[8\] cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__or2_1
Xfanout1001 net1004 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 cpu.SR1.enable vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_8
X_10165_ _05428_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__nand3_1
Xfanout1023 cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_4
Xfanout1034 net1036 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13389__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1045 net1047 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 net1058 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_2
X_10096_ net625 _05131_ net1022 vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__o21a_1
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_2
XANTENNA__14634__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_2
Xfanout1089 net1090 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_2
XANTENNA__09153__B2 _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ clknet_leaf_95_clk _01037_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06767__X _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13855_ clknet_leaf_0_clk _00968_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11325__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ clknet_leaf_38_clk _00025_ net1262 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08982__X _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ a1.CPU_DAT_I\[21\] net928 net276 _05884_ vssd1 vssd1 vccd1 vccd1 _00429_
+ sky130_fd_sc_hd__a22o_1
X_13786_ clknet_leaf_96_clk _00899_ net1231 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ cpu.f0.i\[2\] _06329_ _01872_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XANTENNA__08664__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12668_ net2220 net2126 net1005 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__mux2_1
XANTENNA__06943__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14014__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ clknet_leaf_35_clk _01518_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ net1704 _05817_ net359 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XANTENNA__11015__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ cpu.LCD0.row_2\[1\] net1639 net1012 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XANTENNA__11060__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06662__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12763__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14338_ clknet_leaf_48_clk _01451_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07477__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 cpu.RF0.registers\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10774__A1 cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 cpu.RF0.registers\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 cpu.RF0.registers\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 cpu.RF0.registers\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ clknet_leaf_88_clk _01382_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14164__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09916__B1 cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ _04108_ _04113_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11068__A_N cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1206 cpu.RF0.registers\[9\]\[20\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net300 _03566_ _03538_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__a21oi_1
Xhold1217 cpu.LCD0.row_1\[107\] vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 cpu.LCD0.row_2\[74\] vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 cpu.RF0.registers\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
X_07712_ net956 cpu.RF0.registers\[8\]\[17\] net811 vssd1 vssd1 vccd1 vccd1 _03003_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14231__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ _03980_ _03981_ _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07643_ cpu.RF0.registers\[7\]\[13\] net596 _02908_ _02914_ net624 vssd1 vssd1 vccd1
+ vccd1 _02934_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout169_A _05822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ _02833_ _02864_ net544 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__mux2_2
XFILLER_0_76_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09313_ _03268_ net447 _04243_ _04275_ net465 net453 vssd1 vssd1 vccd1 vccd1 _04604_
+ sky130_fd_sc_hd__mux4_2
X_06525_ cpu.f0.num\[3\] _01793_ _01819_ cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 _01914_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10927__X _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12581__A2_N _06342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_A _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_09244_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06456_ net1705 _01843_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[13\] sky130_fd_sc_hd__xor2_1
XANTENNA__07949__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06853__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08771__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__nor2_1
X_06387_ cpu.f0.num\[12\] vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1245_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14507__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08126_ net1078 cpu.RF0.registers\[28\]\[23\] net867 vssd1 vssd1 vccd1 vccd1 _03417_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10214__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06969__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ net943 cpu.RF0.registers\[10\]\[25\] net860 vssd1 vssd1 vccd1 vccd1 _03348_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09883__B _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__B1 cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ cpu.RF0.registers\[8\]\[23\] net611 _02281_ _02291_ _02296_ vssd1 vssd1 vccd1
+ vccd1 _02299_ sky130_fd_sc_hd__a2111o_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13531__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07933__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09107__C net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net1077 cpu.RF0.registers\[17\]\[26\] net882 vssd1 vssd1 vccd1 vccd1 _04250_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ net1914 net225 net317 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
X_10921_ net2469 net157 net430 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10852_ cpu.DM0.readdata\[7\] net739 net722 vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__o21a_1
X_13640_ clknet_leaf_97_clk _00753_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14037__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10783_ cpu.f0.data_adr\[20\] _05096_ net991 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__mux2_1
X_13571_ clknet_leaf_79_clk _00684_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08110__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ cpu.DM0.dhit _06249_ cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__a21o_1
XANTENNA__13061__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10285__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14187__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11404_ net2515 net249 net384 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12384_ net1119 net1853 net529 cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1 vccd1 _01510_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10756__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10756__B2 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14123_ clknet_leaf_91_clk _01236_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11335_ net503 _05912_ _05920_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__and3_1
XANTENNA__12704__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06975__A3 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ net2538 net138 net402 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__mux2_1
X_14054_ clknet_leaf_8_clk _01167_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08042__X _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ clknet_leaf_36_clk _00194_ net1260 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
X_10217_ net725 _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__and2_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11197_ net1577 net148 net410 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07881__X _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ _05414_ _05415_ cpu.IM0.address_IM\[25\] net1022 vssd1 vssd1 vccd1 vccd1
+ _00048_ sky130_fd_sc_hd__o2bb2a_1
X_10079_ _05346_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__and2_1
XANTENNA__06938__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07137__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_67_clk _01020_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07760__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11055__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ clknet_leaf_1_clk _00951_ net1139 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12433__A1 cpu.DM0.readdata\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ clknet_leaf_104_clk _00882_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_80_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08101__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13404__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10444__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07290_ net545 _02579_ _02580_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_80_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06673__A a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13554__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 cpu.RF0.registers\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 cpu.RF0.registers\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold325 cpu.RF0.registers\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 cpu.RF0.registers\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 cpu.RF0.registers\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold358 cpu.RF0.registers\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _05214_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nor2_1
Xhold369 cpu.RF0.registers\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload23_A clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 _02143_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__A1 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08168__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout816 net819 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
X_09862_ _02719_ _02720_ _01786_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a21o_1
Xfanout827 _02129_ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_4
XFILLER_0_0_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout838 _02052_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_2
Xfanout849 _02041_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_6
Xhold1003 a1.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net938 cpu.RF0.registers\[8\]\[19\] net873 vssd1 vssd1 vccd1 vccd1 _04104_
+ sky130_fd_sc_hd__and3_1
X_09793_ net303 _05083_ _05082_ net277 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a2bb2o_1
Xhold1014 cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 cpu.LCD0.row_1\[59\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 cpu.RF0.registers\[9\]\[28\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 _01685_ vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _04031_ _04032_ _03869_ _03902_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a211o_1
Xhold1058 cpu.RF0.registers\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__A2 _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 cpu.RF0.registers\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ net471 _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07670__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1195_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ net1045 cpu.RF0.registers\[28\]\[13\] net765 vssd1 vssd1 vccd1 vccd1 _02917_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08628__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ cpu.RF0.registers\[5\]\[8\] net602 net579 cpu.RF0.registers\[18\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__a22o_1
XANTENNA__13084__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06508_ cpu.f0.num\[25\] cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07679__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07488_ net1060 cpu.RF0.registers\[19\]\[5\] net823 vssd1 vssd1 vccd1 vccd1 _02779_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07300__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__A1 _02381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06439_ cpu.CU0.opcode\[3\] cpu.CU0.opcode\[2\] cpu.CU0.opcode\[1\] cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__or4bb_4
X_09227_ _03302_ _04289_ _04292_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__A1 cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1150_X net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12188__B1 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07829__D _03119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ _02093_ _02108_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08109_ _03391_ _03392_ _03397_ _03399_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__or4_1
X_09089_ _02099_ _02106_ _02110_ _02112_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__or4_4
XANTENNA__12921__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120_ net1720 net189 net418 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold870 cpu.RF0.registers\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12821__Q cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 cpu.RF0.registers\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net2148 net175 net428 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold892 cpu.RF0.registers\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09118__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ _05259_ _05261_ _05267_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_53_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12112__B1 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11953_ net2771 net153 net318 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__mux2_1
XANTENNA__07580__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08867__B1 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08331__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13427__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10904_ net1550 net169 net430 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
X_14672_ net1394 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_101_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ net2377 net181 net328 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ clknet_leaf_65_clk _00736_ net1282 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ cpu.DM0.readdata\[2\] _05043_ net739 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_24_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11603__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13554_ clknet_leaf_70_clk _00667_ net1326 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10766_ net987 cpu.f0.data_adr\[15\] vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13577__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12505_ _05540_ _06268_ _06285_ net262 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__o211a_1
X_10697_ net2557 net2402 net902 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ clknet_leaf_101_clk _00598_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12179__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12436_ cpu.DM0.data_i\[26\] net534 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08398__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net1120 net1454 net530 cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ clknet_leaf_86_clk _01219_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11318_ net2203 net175 net396 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__mux2_1
X_12298_ net112 net555 vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__or2_1
X_14037_ clknet_leaf_74_clk _01150_ net1324 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11249_ net2908 net197 net402 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14202__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08570__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ _02070_ _02075_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__or3_1
XANTENNA__06668__A a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08586__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09044__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08858__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08460_ cpu.RF0.registers\[4\]\[8\] net678 _03748_ _03749_ _03750_ vssd1 vssd1 vccd1
+ vccd1 _03751_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14352__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07411_ net1048 cpu.RF0.registers\[31\]\[0\] net830 vssd1 vssd1 vccd1 vccd1 _02702_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08391_ cpu.RF0.registers\[8\]\[10\] net708 net691 cpu.RF0.registers\[10\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_15_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11513__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07342_ cpu.RF0.registers\[28\]\[3\] net577 _02613_ _02620_ _02626_ vssd1 vssd1 vccd1
+ vccd1 _02633_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10968__A1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14393__Q cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07273_ net1061 cpu.RF0.registers\[25\]\[7\] net759 vssd1 vssd1 vccd1 vccd1 _02564_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09012_ net1074 cpu.RF0.registers\[18\]\[31\] net855 vssd1 vssd1 vccd1 vccd1 _04303_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12944__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07786__X _03077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold100 _00172_ vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09586__A1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold111 _00153_ vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _00183_ vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06850__B net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 cpu.f0.write_data\[26\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__B1 _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 cpu.RF0.registers\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 cpu.f0.read_i vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07665__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold166 cpu.RF0.registers\[0\]\[6\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _00336_ vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold188 a1.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 a1.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _05149_ _05198_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a21oi_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_8
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_8
Xfanout624 _02127_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1110_A cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net637 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout646 _02061_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ net298 _04945_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__nand2_1
Xfanout657 _02054_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout570_A _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _02050_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
Xfanout679 _02037_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A _02050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _02795_ net436 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__nor2_1
X_06988_ net1034 cpu.RF0.registers\[31\]\[23\] net825 vssd1 vssd1 vccd1 vccd1 _02279_
+ sky130_fd_sc_hd__and3_1
X_08727_ cpu.RF0.registers\[12\]\[0\] net946 net868 vssd1 vssd1 vccd1 vccd1 _04018_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09889__A cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ net1102 cpu.RF0.registers\[21\]\[2\] _02019_ vssd1 vssd1 vccd1 vccd1 _03949_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10120__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09241__X _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07609_ _02895_ _02896_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08589_ net949 cpu.RF0.registers\[12\]\[4\] net868 vssd1 vssd1 vccd1 vccd1 _03880_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11423__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ net2263 cpu.LCD0.row_1\[34\] net897 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10959__A1 _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12816__Q cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ net52 net921 vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10482_ net98 net923 net748 net1513 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__a22o_1
X_13270_ clknet_leaf_23_clk cpu.RU0.next_FetchedInstr\[9\] net1178 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_92_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12221_ cpu.LCD0.row_1\[68\] _06001_ _06012_ cpu.LCD0.row_2\[108\] _06117_ vssd1
+ vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_92_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06760__B net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ cpu.LCD0.row_2\[97\] _06018_ _06034_ cpu.LCD0.row_2\[25\] vssd1 vssd1 vccd1
+ vccd1 _06052_ sky130_fd_sc_hd__a22o_1
XANTENNA__07052__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14225__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ net2048 net237 net420 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12083_ _01773_ cpu.LCD0.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__nor2_2
XANTENNA__08968__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11034_ cpu.IG0.Instr\[8\] cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__and2b_2
XFILLER_0_60_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12833__SET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14375__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ clknet_leaf_28_clk _00174_ net1188 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09501__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ net1807 net229 net320 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XANTENNA__06775__X _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09151__X _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14655_ clknet_leaf_61_clk _01756_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ net2862 net248 net328 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__mux2_1
XANTENNA__12967__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11333__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ clknet_leaf_7_clk _00719_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10818_ cpu.IM0.address_IM\[30\] net1013 net284 _05759_ vssd1 vssd1 vccd1 vccd1 _05760_
+ sky130_fd_sc_hd__a22o_1
X_14586_ clknet_leaf_51_clk _01688_ net1377 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_11798_ net2786 net236 net336 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13537_ clknet_leaf_63_clk _00650_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10749_ net287 _05709_ _05710_ net1016 cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1
+ vccd1 _05711_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07469__D _02756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09017__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07291__A2 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ clknet_leaf_8_clk _00581_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12851__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ net2463 net730 net500 _06233_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__o22a_1
XANTENNA__06670__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13399_ clknet_leaf_65_clk _00512_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07485__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ net1098 cpu.RF0.registers\[18\]\[29\] net853 vssd1 vssd1 vccd1 vccd1 _03251_
+ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_4_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08878__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__X _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ cpu.RF0.registers\[4\]\[27\] net586 _02188_ _02156_ _02163_ vssd1 vssd1 vccd1
+ vccd1 _02202_ sky130_fd_sc_hd__a2111o_1
X_07891_ cpu.RF0.registers\[26\]\[29\] net600 _02191_ cpu.RF0.registers\[25\]\[29\]
+ _03175_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11508__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14667__1389 vssd1 vssd1 vccd1 vccd1 _14667__1389/HI net1389 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_88_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09630_ _04647_ _04915_ _04918_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__or4_1
X_06842_ net1038 cpu.RF0.registers\[19\]\[27\] net821 vssd1 vssd1 vccd1 vccd1 _02133_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ net294 _04849_ _04850_ net297 _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__o221a_1
X_06773_ net1084 net836 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_65_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08512_ _03797_ _03800_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__and2_1
X_09492_ _04781_ _04782_ net475 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload90_A clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07503__B1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08443_ _03729_ _03731_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout151_A _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _05774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11243__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _02832_ _02867_ net491 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13892__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07325_ net974 cpu.RF0.registers\[2\]\[3\] net772 vssd1 vssd1 vccd1 vccd1 _02616_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1060_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10810__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07256_ net1062 cpu.RF0.registers\[30\]\[7\] net763 vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07282__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14248__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07187_ net1046 cpu.RF0.registers\[25\]\[10\] net757 vssd1 vssd1 vccd1 vccd1 _02478_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_83_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10169__A2 _04601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08782__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13272__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14398__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout410 _05917_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
Xfanout421 _05914_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
XANTENNA__07692__A _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_6
Xfanout443 _03505_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout454 _02756_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net469 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_4
XANTENNA__08534__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ _04753_ _04813_ _04830_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__nand3_1
Xfanout487 _02642_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_2
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07742__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _05044_ _05046_ _05049_ net304 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ cpu.f0.write_data\[28\] net498 net279 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1
+ _01749_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ net2167 net164 net346 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11153__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ clknet_leaf_28_clk _01550_ net1188 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11652_ net1493 net171 net355 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ net2130 cpu.LCD0.row_1\[17\] net908 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ clknet_leaf_26_clk _01482_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11583_ net1743 net205 net362 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13322_ clknet_leaf_23_clk cpu.RU0.next_FetchedData\[29\] net1178 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[29\] sky130_fd_sc_hd__dfrtp_1
X_10534_ net1133 net1613 net913 _05654_ vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_2
X_13253_ clknet_leaf_36_clk _00433_ net1263 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ net15 net754 net564 net1825 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a22o_1
X_12204_ _06085_ _06087_ _06089_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ clknet_leaf_36_clk _00364_ net1265 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ net1126 _01801_ net266 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12135_ net745 _05981_ _05993_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12712__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ cpu.LCD0.cnt_500hz\[10\] _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__or2_1
XANTENNA__11328__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net2077 net925 net273 _05897_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__a22o_1
XANTENNA__07733__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__A1 cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ clknet_leaf_44_clk net1474 net1305 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10096__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net2045 net164 net322 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06665__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ clknet_leaf_26_clk _00088_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11063__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07500__A3 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14638_ clknet_leaf_24_clk _01739_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13145__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11998__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14569_ clknet_leaf_50_clk _01671_ net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10399__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ net1049 cpu.RF0.registers\[31\]\[14\] net829 net575 cpu.RF0.registers\[14\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_77_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ net938 cpu.RF0.registers\[11\]\[22\] net880 vssd1 vssd1 vccd1 vccd1 _03381_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload20 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__10915__B _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07041_ net1040 cpu.RF0.registers\[16\]\[19\] net831 vssd1 vssd1 vccd1 vccd1 _02332_
+ sky130_fd_sc_hd__and3_1
Xclkload31 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__13295__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload42 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload53 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload53/X sky130_fd_sc_hd__clkbuf_4
Xclkload64 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__14540__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload75 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__inv_6
XANTENNA__07016__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload86 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_3_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload97 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_8
X_08992_ _04275_ _04277_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__or2_1
XANTENNA__07972__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__inv_2
XANTENNA__10859__A0 _05229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A1 _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ cpu.RF0.registers\[3\]\[28\] net609 net602 cpu.RF0.registers\[5\]\[28\] _03164_
+ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09613_ _04710_ _04903_ _04902_ _04897_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__o211a_1
X_06825_ cpu.CU0.funct3\[1\] _02104_ _02107_ _02093_ _02114_ vssd1 vssd1 vccd1 vccd1
+ _02116_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout366_A _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ _04761_ _04834_ net472 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux2_1
X_06756_ net1075 net851 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09232__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__A1 cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ net442 net295 _04402_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a21oi_1
X_06687_ net1712 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[23\] sky130_fd_sc_hd__and2_1
XANTENNA__10378__A cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1275_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__Y _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08426_ cpu.RF0.registers\[9\]\[9\] net699 net648 cpu.RF0.registers\[25\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09229__A0 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ cpu.RF0.registers\[30\]\[11\] net660 net646 cpu.RF0.registers\[21\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_6
XANTENNA__13638__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07308_ cpu.RF0.registers\[23\]\[4\] net613 net587 cpu.RF0.registers\[4\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ cpu.RF0.registers\[10\]\[13\] net691 net654 cpu.RF0.registers\[2\]\[13\]
+ _03575_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a221o_1
XANTENNA__10825__B cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07239_ net1036 cpu.RF0.registers\[28\]\[9\] net765 vssd1 vssd1 vccd1 vccd1 _02530_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10250_ cpu.f0.i\[11\] net541 vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13788__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ net126 _05445_ _05442_ net631 vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a211o_1
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07963__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1216 net1219 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08311__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1227 net1228 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
Xfanout1238 net1241 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13018__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1249 net1255 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _05774_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11148__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 _06252_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout273 _05846_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
X_13940_ clknet_leaf_71_clk _01053_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout284 _05688_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10314__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _04396_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10987__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_87_clk _00984_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09468__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ clknet_leaf_41_clk _00041_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12120__X _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__A1 _05328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14413__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ net1489 net497 net280 cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08140__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11704_ net2015 net234 net347 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
X_12684_ net2760 net2605 net1005 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XANTENNA__07494__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14423_ clknet_leaf_17_clk _01534_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_11635_ net1961 net249 net356 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11578__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07597__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14563__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14354_ clknet_leaf_58_clk _01467_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14666__1388 vssd1 vssd1 vccd1 vccd1 _14666__1388/HI net1388 sky130_fd_sc_hd__conb_1
X_11566_ net505 _05907_ _05910_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__and3_4
XFILLER_0_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14491__Q cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13305_ clknet_leaf_31_clk cpu.RU0.next_FetchedData\[12\] net1205 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06932__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ net65 net917 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__and2_1
XANTENNA__10227__S net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14285_ clknet_leaf_103_clk _01398_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11497_ net1947 net140 net376 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13236_ clknet_leaf_43_clk _00416_ net1303 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10448_ net28 net753 net563 a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09943__A1 cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ clknet_leaf_37_clk _00347_ net1260 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ net1126 _05607_ net266 net1889 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12118_ net745 _05984_ _05987_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__and3_4
XANTENNA__09317__A _03119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ clknet_leaf_52_clk _00278_ net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07763__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11058__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12049_ _01956_ _05957_ _05961_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__and3_1
XANTENNA__10897__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06610_ _01974_ _01755_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__xnor2_1
X_07590_ net968 cpu.RF0.registers\[11\]\[12\] net779 vssd1 vssd1 vccd1 vccd1 _02881_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06676__A a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14093__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06541_ _01926_ _01927_ _01928_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06472_ _01780_ _01791_ vssd1 vssd1 vccd1 vccd1 cpu.DM0.next_enable sky130_fd_sc_hd__nor2_2
XANTENNA__09987__A cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ net493 _04518_ _04519_ _04550_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11018__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ cpu.RF0.registers\[22\]\[21\] net670 net666 _03489_ _03501_ vssd1 vssd1 vccd1
+ vccd1 _03502_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09191_ net303 _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07003__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11521__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ _03420_ _03421_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__nor4_1
XANTENNA__08434__A1 cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__A2 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload53_A clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06842__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ _03360_ _03361_ _03362_ _03363_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__or4_1
XANTENNA__13930__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07024_ net1086 _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10544__A2 a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1023_A cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ cpu.RF0.registers\[20\]\[26\] net710 net654 cpu.RF0.registers\[2\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a22o_1
XANTENNA__07673__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 cpu.RF0.registers\[0\]\[12\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _01717_ vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 cpu.f0.data_adr\[21\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ net1030 cpu.RF0.registers\[31\]\[30\] net826 vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__and3_1
Xhold48 cpu.FetchedInstr\[9\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 _00154_ vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14436__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _02274_ _02312_ net259 _03145_ net488 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__A cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08370__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ _02094_ _02098_ _02092_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06920__A1 cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ _03077_ _03078_ net522 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09527_ _02508_ net435 net289 _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06739_ net1087 net859 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__and2_2
XANTENNA__14178__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_X net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13460__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14586__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__A cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _04747_ _04748_ _04745_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14107__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A1 cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11009__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ _02508_ _03665_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__xnor2_1
X_09389_ _04597_ _04671_ net481 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ net2124 net187 net384 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XANTENNA__12221__A2 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_X clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__A _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__Q cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ net2845 net173 net392 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10302_ net1020 _05539_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__and2_1
X_14070_ clknet_leaf_59_clk _01183_ net1348 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11282_ net1771 net208 net399 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__mux2_1
XANTENNA__13742__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ clknet_leaf_34_clk _00210_ net1253 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
X_10233_ cpu.f0.i\[8\] cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__nand2_1
XANTENNA__12115__X _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08679__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ cpu.IM0.address_IM\[26\] _02248_ _05419_ vssd1 vssd1 vccd1 vccd1 _05430_
+ sky130_fd_sc_hd__a21o_1
Xfanout1013 net1017 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07583__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1024 net1025 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_2
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_2
XFILLER_0_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_41_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10095_ net125 _05364_ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a21o_1
XANTENNA__12288__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 cpu.IG0.Instr\[22\] vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_4
Xfanout1079 net1091 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_2
X_13923_ clknet_leaf_78_clk _01036_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08361__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08900__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13854_ clknet_leaf_85_clk _00967_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13803__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14486__Q cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ net2834 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_28_clk_X clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13785_ clknet_leaf_92_clk _00898_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10997_ cpu.f0.write_data\[21\] _05883_ net993 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__mux2_1
X_12736_ _06326_ _01762_ _01765_ net498 cpu.f0.write_data\[1\] vssd1 vssd1 vccd1 vccd1
+ _01722_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_100_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ cpu.LCD0.row_2\[69\] cpu.LCD0.row_2\[61\] net997 vssd1 vssd1 vccd1 vccd1
+ _01660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07872__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ clknet_leaf_35_clk _01517_ net1258 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ net2423 net187 net360 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
X_12598_ cpu.LCD0.row_2\[0\] net1641 net1012 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XANTENNA__07758__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14337_ clknet_leaf_48_clk _01450_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10223__B2 cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11549_ net2081 net175 net368 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14309__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 a1.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10774__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold518 cpu.RF0.registers\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 cpu.RF0.registers\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ clknet_leaf_14_clk _01381_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap259 _03120_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_1
XANTENNA__08719__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13219_ clknet_leaf_6_clk _00399_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09916__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14199_ clknet_leaf_65_clk _01312_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08589__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14459__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13333__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1207 cpu.RF0.registers\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _03802_ _04039_ _04047_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a31o_2
XANTENNA__12279__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1218 _00323_ vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1229 _01665_ vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07711_ net1027 cpu.RF0.registers\[22\]\[17\] net799 vssd1 vssd1 vccd1 vccd1 _03002_
+ sky130_fd_sc_hd__and3_1
X_08691_ cpu.RF0.registers\[5\]\[1\] net704 _02033_ cpu.RF0.registers\[15\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11516__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07642_ _02929_ _02930_ _02931_ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ _02861_ _02862_ _02863_ net619 cpu.RF0.registers\[0\]\[8\] vssd1 vssd1 vccd1
+ vccd1 _02864_ sky130_fd_sc_hd__o32a_2
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08104__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09447__A3 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ net446 _03371_ _03402_ net445 net460 net454 vssd1 vssd1 vccd1 vccd1 _04603_
+ sky130_fd_sc_hd__mux4_2
X_06524_ cpu.f0.num\[5\] _01795_ cpu.f0.num\[10\] _01801_ _01912_ vssd1 vssd1 vccd1
+ vccd1 _01913_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07458__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09510__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__A1_N net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ net462 _03992_ _04026_ net456 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o211a_1
X_06455_ _01843_ _01857_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[12\] sky130_fd_sc_hd__nor2_1
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout231_A _05783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06853__B net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__A1 cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06386_ cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__inv_2
X_09174_ net463 _03899_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__nor2_1
XANTENNA__12203__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07668__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07030__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10214__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08125_ net935 cpu.RF0.registers\[9\]\[23\] net862 vssd1 vssd1 vccd1 vccd1 _03416_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ net1087 cpu.RF0.registers\[21\]\[25\] net865 vssd1 vssd1 vccd1 vccd1 _03347_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09368__C1 _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ net1034 cpu.RF0.registers\[30\]\[23\] net761 vssd1 vssd1 vccd1 vccd1 _02298_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09907__B2 cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_40_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A _02019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net936 cpu.RF0.registers\[1\]\[26\] net882 vssd1 vssd1 vccd1 vccd1 _04249_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13826__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ net957 cpu.RF0.registers\[6\]\[30\] net800 vssd1 vssd1 vccd1 vccd1 _03200_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ cpu.RF0.registers\[28\]\[17\] net705 net642 cpu.RF0.registers\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11426__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _05424_ _05833_ net719 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12850__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12819__Q cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ net740 _04880_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ clknet_leaf_102_clk _00683_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10782_ a1.ADR_I\[19\] net560 net538 _05734_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09420__A _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ cpu.f0.i\[25\] _06294_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_40_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13206__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11161__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12452_ net1129 cpu.f0.state\[3\] _06249_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_87_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10205__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08949__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ net2925 net256 net385 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10853__X _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12383_ net1119 net2652 net529 cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 _01509_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14122_ clknet_leaf_100_clk _01235_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09419__X _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ cpu.RF0.registers\[9\]\[31\] net129 net394 vssd1 vssd1 vccd1 vccd1 _00759_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13356__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14601__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ clknet_leaf_3_clk _01166_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11265_ net2260 net140 net404 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
XANTENNA__10508__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ clknet_leaf_36_clk _00193_ net1263 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
X_10216_ net527 net307 vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__or2_1
X_11196_ net2609 net155 net410 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__mux2_1
XANTENNA__08582__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12720__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ net625 _04663_ net1022 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09126__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _05328_ _05348_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11336__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13906_ clknet_leaf_61_clk _01019_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07688__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ clknet_leaf_103_clk _00950_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09033__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13768_ clknet_leaf_97_clk _00881_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10444__B2 a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12719_ net1491 cpu.LCD0.row_2\[113\] net1011 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ clknet_leaf_78_clk _00812_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06673__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11071__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14131__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07860__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 cpu.DM0.readdata\[3\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07612__A2 _02901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 cpu.RF0.registers\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14281__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold326 cpu.RF0.registers\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 cpu.RF0.registers\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 cpu.RF0.registers\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _05205_ _05206_ _05204_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold359 cpu.RF0.registers\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13849__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net809 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
XANTENNA_wire833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09861_ _02719_ _02720_ _01786_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a21oi_1
Xfanout817 net819 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_4
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload16_A clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 _02052_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_8
X_08812_ cpu.RF0.registers\[2\]\[19\] net654 _04100_ _04101_ _04102_ vssd1 vssd1 vccd1
+ vccd1 _04103_ sky130_fd_sc_hd__a2111o_1
X_09792_ _04413_ _04488_ _04489_ net292 _04770_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1004 cpu.RF0.registers\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 cpu.RF0.registers\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1026 cpu.RF0.registers\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ _04031_ _04032_ _03902_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a21o_1
XANTENNA__12873__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 cpu.RF0.registers\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07951__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1048 cpu.RF0.registers\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 cpu.LCD0.row_2\[23\] vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06848__B net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08674_ net468 net458 net492 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__a21oi_1
X_07625_ net964 cpu.RF0.registers\[6\]\[13\] net800 vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10938__X _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07556_ net973 cpu.RF0.registers\[13\]\[8\] net793 vssd1 vssd1 vccd1 vccd1 _02847_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06864__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ cpu.f0.num\[16\] cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10386__A cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ net982 cpu.RF0.registers\[15\]\[5\] net828 vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1355_A net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09226_ net511 _04294_ _04453_ _04515_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o31ai_4
X_06438_ cpu.CU0.opcode\[2\] cpu.CU0.opcode\[0\] cpu.CU0.opcode\[1\] vssd1 vssd1 vccd1
+ vccd1 _01846_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13379__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14624__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09157_ net511 _04363_ _04364_ _04445_ cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1
+ _04448_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_20_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06369_ cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1143_X net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07695__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ cpu.RF0.registers\[16\]\[22\] net636 _03386_ _03398_ net665 vssd1 vssd1 vccd1
+ vccd1 _03399_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_82_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09088_ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__inv_2
XANTENNA__08143__X _03434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06811__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ cpu.RF0.registers\[8\]\[24\] _02014_ net644 cpu.RF0.registers\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 cpu.LCD0.row_2\[110\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 cpu.LCD0.row_1\[23\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold882 cpu.LCD0.row_1\[17\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold893 cpu.LCD0.row_2\[54\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net2666 net196 net428 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ cpu.IM0.address_IM\[13\] _02904_ _05279_ vssd1 vssd1 vccd1 vccd1 _05280_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08022__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07906__A3 _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14004__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11156__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ net2744 net163 net318 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__mux2_1
XANTENNA__08867__A1 cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ net722 _05365_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__o21ai_4
X_14671_ net1393 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_11883_ net1679 net172 net327 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14154__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ clknet_leaf_58_clk _00735_ net1368 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net2034 net253 net431 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XANTENNA__06774__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12415__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ clknet_leaf_76_clk _00666_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ net990 _05140_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__nand2_1
XANTENNA__08095__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10977__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _05540_ _06268_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nor2_1
XANTENNA__07842__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13484_ clknet_leaf_80_clk _00597_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10696_ cpu.LCD0.row_1\[102\] net2429 net908 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12435_ net2616 net730 net500 _06241_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09149__X _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12366_ net1119 net1733 net529 cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 _01492_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06940__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14105_ clknet_leaf_92_clk _01218_ net1240 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11317_ net2302 net194 net396 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12297_ _06173_ _06175_ _06177_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__or4_2
X_14036_ clknet_leaf_73_clk _01149_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12896__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ net2432 net208 net403 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__mux2_1
X_11179_ cpu.RF0.registers\[5\]\[9\] net216 net410 vssd1 vssd1 vccd1 vccd1 _00609_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07771__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06668__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07410_ net1048 cpu.RF0.registers\[22\]\[0\] net803 vssd1 vssd1 vccd1 vccd1 _02701_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09807__A0 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ net1093 cpu.RF0.registers\[31\]\[10\] net857 vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13521__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07341_ cpu.RF0.registers\[18\]\[3\] net579 _02619_ _02623_ _02630_ vssd1 vssd1 vccd1
+ vccd1 _02632_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14647__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07272_ net1062 cpu.RF0.registers\[19\]\[7\] net823 vssd1 vssd1 vccd1 vccd1 _02563_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07833__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09011_ net934 cpu.RF0.registers\[7\]\[31\] net844 vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 cpu.LCD0.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 net104 vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 cpu.LCD0.row_2\[127\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold134 cpu.RF0.registers\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold145 cpu.RF0.registers\[0\]\[5\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 a1.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold167 cpu.RF0.registers\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net717 net134 _05199_ net631 vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a31o_1
Xhold178 cpu.LCD0.row_2\[26\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _02148_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_8
XANTENNA__14027__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 cpu.RF0.registers\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout614 _02135_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_8
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_A _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout636 _02066_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_6
X_09844_ _04411_ _04697_ _05134_ net305 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__o22a_1
Xfanout647 _02061_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
Xfanout658 _02054_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10353__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07307__X _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__C _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ _05063_ _05065_ net306 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06987_ net955 cpu.RF0.registers\[5\]\[23\] net795 vssd1 vssd1 vccd1 vccd1 _02278_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13051__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ cpu.RF0.registers\[5\]\[0\] net703 _04014_ _04015_ _04016_ vssd1 vssd1 vccd1
+ vccd1 _04017_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09522__X _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ net1102 cpu.RF0.registers\[28\]\[2\] net868 vssd1 vssd1 vccd1 vccd1 _03948_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09889__B cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ cpu.RF0.registers\[17\]\[12\] net605 _02870_ _02898_ net621 vssd1 vssd1 vccd1
+ vccd1 _02899_ sky130_fd_sc_hd__a2111o_1
X_08588_ net1101 cpu.RF0.registers\[27\]\[4\] net879 vssd1 vssd1 vccd1 vccd1 _03879_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10828__B _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07539_ _02797_ _02829_ net545 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__mux2_4
XFILLER_0_7_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10959__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ net1133 a1.ADR_I\[19\] net913 _05662_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07824__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08017__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09209_ _04498_ _04499_ net454 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__mux2_1
X_10481_ net1464 net923 net748 a1.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22o_1
XANTENNA__10844__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12220_ cpu.LCD0.row_1\[84\] _05986_ _06033_ cpu.LCD0.row_2\[76\] vssd1 vssd1 vccd1
+ vccd1 _06117_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10563__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12832__Q cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12581__B2 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ cpu.LCD0.row_2\[57\] _06000_ _06049_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09129__B _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__B1 _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ _05765_ _05907_ net503 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and3_4
X_12082_ net746 _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__and3_4
Xhold690 cpu.RF0.registers\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _05763_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__and2_1
XANTENNA__12123__X _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14303__RESET_B net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06769__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__X _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ clknet_leaf_44_clk net1486 net1305 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
Xhold1390 cpu.RF0.registers\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13544__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11935_ net1676 net232 net320 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14654_ clknet_leaf_61_clk _01755_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11866_ net1686 net252 net328 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14494__Q cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06935__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ clknet_leaf_2_clk _00718_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ cpu.f0.data_adr\[30\] _04517_ net989 vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__mux2_1
X_14585_ clknet_leaf_50_clk _01687_ net1384 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11797_ net506 _05906_ _05920_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and3_4
XFILLER_0_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13536_ clknet_leaf_9_clk _00649_ net1160 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10748_ net992 cpu.f0.data_adr\[10\] vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07815__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13467_ clknet_leaf_92_clk _00580_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10679_ cpu.LCD0.row_1\[85\] cpu.LCD0.row_1\[93\] net900 vssd1 vssd1 vccd1 vccd1
+ _00309_ sky130_fd_sc_hd__mux2_1
XANTENNA__10754__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07539__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__X _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ cpu.DM0.data_i\[17\] net534 vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07766__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ clknet_leaf_71_clk _00511_ net1340 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ cpu.LCD0.cnt_20ms\[16\] cpu.LCD0.cnt_20ms\[15\] _06213_ vssd1 vssd1 vccd1
+ vccd1 _06217_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08240__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13074__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ cpu.RF0.registers\[17\]\[27\] net605 _02161_ _02180_ _02133_ vssd1 vssd1
+ vccd1 vccd1 _02201_ sky130_fd_sc_hd__a2111o_1
X_14019_ clknet_leaf_78_clk _01132_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_07890_ cpu.RF0.registers\[27\]\[29\] net592 net571 cpu.RF0.registers\[12\]\[29\]
+ _03178_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__a221o_1
XANTENNA__06679__A a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09055__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ net1042 net822 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__and2_1
XANTENNA__10886__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__A1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09560_ _04391_ _04405_ _04848_ net435 _02866_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_84_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06772_ net944 _02062_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09491_ _04719_ _04759_ net456 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__mux2_1
XANTENNA__07503__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07006__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11524__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08700__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ _03729_ _03731_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nor2_1
XANTENNA__12911__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload83_A clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06845__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ cpu.IM0.address_IM\[11\] net552 _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_
+ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_22_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout144_A _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07324_ net975 cpu.RF0.registers\[14\]\[3\] net763 vssd1 vssd1 vccd1 vccd1 _02615_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12260__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07255_ net1061 cpu.RF0.registers\[28\]\[7\] net767 vssd1 vssd1 vccd1 vccd1 _02546_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout311_A _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07019__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ net1051 cpu.RF0.registers\[26\]\[10\] net787 vssd1 vssd1 vccd1 vccd1 _02477_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13417__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1220_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08231__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1318_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout680_A _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout400 _05921_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout411 _05917_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout422 net425 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _05767_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
Xfanout444 _03471_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
Xfanout477 _02680_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_2
XANTENNA__10877__A1 _05086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _04792_ _05086_ _05107_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__or4_1
XANTENNA__13567__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout488 net490 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
Xfanout499 _01761_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _04384_ _05047_ _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06876__X _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08709_ cpu.RF0.registers\[9\]\[0\] net700 net695 cpu.RF0.registers\[17\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _03833_ _02830_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ net1879 net167 net349 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08309__A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06755__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12827__Q cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11651_ net2766 net187 net357 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ net2457 cpu.LCD0.row_1\[16\] net909 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
X_14370_ clknet_leaf_27_clk cpu.K0.next_keyvalid net1183 vssd1 vssd1 vccd1 vccd1 cpu.K0.keyvalid
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12251__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ net2096 net175 net364 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ clknet_leaf_17_clk cpu.RU0.next_FetchedData\[28\] net1195 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[28\] sky130_fd_sc_hd__dfrtp_1
X_10533_ net42 net920 vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12118__X _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire856 _02035_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_44_clk _00432_ net1305 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06481__A1 cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire878 _02010_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_2
X_10464_ net14 net752 net562 net1422 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__o22a_1
XANTENNA__07586__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13097__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12203_ cpu.LCD0.row_1\[123\] _06014_ _06091_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_
+ sky130_fd_sc_hd__a211o_1
X_13183_ clknet_leaf_34_clk _00363_ net1253 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ net1125 _05615_ net264 net2732 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__a2bb2o_1
X_12134_ cpu.LCD0.row_2\[72\] _06033_ _06034_ cpu.LCD0.row_2\[24\] vssd1 vssd1 vccd1
+ vccd1 _06035_ sky130_fd_sc_hd__a22o_1
XANTENNA__11609__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12065_ _05971_ net502 _05970_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__and3b_1
XFILLER_0_25_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14489__Q cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ cpu.f0.write_data\[27\] _05896_ net985 vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__mux2_1
XANTENNA__14492__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12967_ clknet_leaf_44_clk net1524 net1312 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08289__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ net2683 net168 net325 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XANTENNA__11293__A1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10096__A2 _05131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ clknet_leaf_27_clk _00087_ net1188 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09041__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11849_ net1844 net185 net332 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
X_14637_ clknet_leaf_21_clk _01738_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14568_ clknet_leaf_46_clk _01670_ net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09789__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08506__X _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08880__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13519_ clknet_leaf_82_clk _00632_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14499_ clknet_leaf_54_clk _01601_ net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload10 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07040_ net963 cpu.RF0.registers\[15\]\[19\] net827 vssd1 vssd1 vccd1 vccd1 _02331_
+ sky130_fd_sc_hd__and3_1
Xclkload21 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload21/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload32 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload32/X sky130_fd_sc_hd__clkbuf_8
Xclkload43 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_4
Xclkload54 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__inv_6
XFILLER_0_80_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload65 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_45_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload76 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08213__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload87 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_8
XFILLER_0_45_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload98 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_12
XFILLER_0_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07793__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ _03371_ _03373_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__o21a_1
XANTENNA__11519__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ net509 _03231_ net522 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14399__Q cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07873_ cpu.RF0.registers\[15\]\[28\] net590 net583 cpu.RF0.registers\[6\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a22o_1
XANTENNA__06527__A2 _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ net472 net272 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nand2_1
XANTENNA__08120__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06824_ net1118 net633 _02113_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09513__A _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _04780_ _04833_ net456 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__mux2_1
X_06755_ net1080 cpu.RF0.registers\[23\]\[30\] net844 vssd1 vssd1 vccd1 vccd1 _02046_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout359_A _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10087__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _02941_ net442 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__nor2_1
X_06686_ net2073 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14215__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07033__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ cpu.RF0.registers\[17\]\[9\] net694 _03701_ _03706_ _03713_ vssd1 vssd1 vccd1
+ vccd1 _03716_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09229__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1268_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08356_ net1088 cpu.RF0.registers\[23\]\[11\] net847 vssd1 vssd1 vccd1 vccd1 _03647_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_12
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07307_ _02591_ _02593_ _02595_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__or4_2
XFILLER_0_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ net937 cpu.RF0.registers\[1\]\[13\] net882 vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10795__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06591__B _01965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14365__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07238_ net1035 cpu.RF0.registers\[23\]\[9\] net816 vssd1 vssd1 vccd1 vccd1 _02529_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09937__C1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08204__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07169_ cpu.RF0.registers\[12\]\[11\] net571 _02441_ _02447_ _02457_ vssd1 vssd1
+ vccd1 vccd1 _02460_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08799__A net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1210 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
Xfanout1217 net1219 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_2
XANTENNA__12957__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout1228 net1268 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net244 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XANTENNA__13948__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1239 net1241 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
Xfanout252 _05774_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout263 _06252_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 net276 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout285 net287 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07176__C1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ clknet_leaf_5_clk _00983_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08965__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ clknet_leaf_15_clk _00040_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09468__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__B net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ net1445 _01761_ net280 cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__X _05001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ net2681 net243 net347 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12683_ cpu.LCD0.row_2\[85\] cpu.LCD0.row_2\[77\] net998 vssd1 vssd1 vccd1 vccd1
+ _01676_ sky130_fd_sc_hd__mux2_1
XANTENNA__10856__X _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08691__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11027__A1 _04357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14422_ clknet_leaf_17_clk _01533_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12224__B1 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ net2143 net253 net356 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08979__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14353_ clknet_leaf_57_clk _01466_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11565_ net2506 net129 net366 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ clknet_leaf_24_clk cpu.RU0.next_FetchedData\[11\] net1204 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[11\] sky130_fd_sc_hd__dfrtp_1
X_10516_ net1134 net1833 net912 _05645_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14284_ clknet_leaf_68_clk _01397_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11496_ net2714 net144 net376 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__mux2_1
XANTENNA__13732__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ clknet_leaf_44_clk _00415_ net1306 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net27 net754 net564 a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ clknet_leaf_35_clk _00346_ net1260 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ cpu.f0.i\[1\] net270 vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__nand2_1
XANTENNA__11339__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ net746 _05981_ net557 vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__and3_4
XFILLER_0_23_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13097_ clknet_leaf_48_clk _00277_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09317__B _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13882__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09156__B1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ cpu.LCD0.cnt_500hz\[0\] cpu.LCD0.cnt_500hz\[1\] cpu.LCD0.cnt_500hz\[2\] cpu.LCD0.cnt_500hz\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__a31o_1
XANTENNA__09036__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08903__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07182__A2 _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ clknet_leaf_87_clk _01112_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11074__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06540_ cpu.f0.num\[9\] _01799_ cpu.f0.num\[11\] _01803_ _01915_ vssd1 vssd1 vccd1
+ vccd1 _01929_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09620__X _04911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06471_ _01865_ _01866_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13262__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ cpu.RF0.registers\[17\]\[21\] net694 net677 cpu.RF0.registers\[4\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11802__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14388__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__A1 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09190_ net485 net437 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07890__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06692__A a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12766__A1 cpu.f0.write_data\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12766__B2 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08141_ cpu.RF0.registers\[15\]\[23\] net682 net654 cpu.RF0.registers\[2\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08434__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ cpu.RF0.registers\[16\]\[25\] net636 _03344_ _03352_ _03353_ vssd1 vssd1
+ vccd1 vccd1 _03363_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07023_ net716 _02085_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09067__X _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A1_N _03469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12930__Q a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ cpu.RF0.registers\[15\]\[26\] net682 net636 cpu.RF0.registers\[16\]\[26\]
+ _04252_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 a1.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 net122 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ net1029 cpu.RF0.registers\[20\]\[30\] net780 vssd1 vssd1 vccd1 vccd1 _03216_
+ sky130_fd_sc_hd__and3_1
Xhold38 cpu.RF0.registers\[0\]\[13\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 cpu.FetchedInstr\[17\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A1 _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _02312_ net259 _03145_ net489 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12588__B _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__X _02606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ cpu.CU0.opcode\[3\] cpu.CU0.funct3\[2\] _02092_ _02096_ vssd1 vssd1 vccd1
+ vccd1 _02098_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07787_ net1071 net633 net519 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout643_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1385_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net294 net296 _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__mux2_1
XANTENNA__11257__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13605__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06738_ net1114 net1116 net1110 net1112 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__and4_4
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09457_ _02983_ net435 _04746_ net294 net288 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o221a_1
X_06669_ a1.CPU_DAT_O\[5\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[5\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09897__B cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__A1 _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__inv_2
XANTENNA__11009__A1 _02271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07881__A0 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _04564_ _04590_ _04593_ _04566_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12757__A1 cpu.f0.write_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13755__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__inv_2
XANTENNA__08425__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10232__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ net2243 net193 net392 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10301_ net1462 net727 _05543_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__o21a_1
XANTENNA__08025__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ net1812 net202 net399 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ clknet_leaf_36_clk _00209_ net1264 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
X_10232_ net1419 net727 _05484_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__Q cpu.f0.data_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
X_10163_ cpu.IM0.address_IM\[27\] _02211_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__or2_1
XANTENNA__09137__B _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1014 net1016 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13135__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input37_A gpio_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_2
X_10094_ net717 net134 _05365_ net630 vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a31o_1
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
X_13922_ clknet_leaf_94_clk _01035_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13853_ clknet_leaf_67_clk _00966_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06911__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13285__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ net2836 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14530__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ _03077_ net533 net283 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__o21ba_1
X_13784_ clknet_leaf_7_clk _00897_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08992__A _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12735_ cpu.f0.i\[1\] _01872_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08664__A2 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11622__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ cpu.LCD0.row_2\[68\] cpu.LCD0.row_2\[60\] net1002 vssd1 vssd1 vccd1 vccd1
+ _01659_ sky130_fd_sc_hd__mux2_1
XANTENNA__09600__B _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12748__A1 cpu.f0.write_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06943__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ clknet_leaf_35_clk _01516_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11617_ cpu.RF0.registers\[18\]\[17\] net192 net358 vssd1 vssd1 vccd1 vccd1 _01033_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09613__A1 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ _01968_ _01993_ _06354_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10223__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ net2479 net196 net368 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
X_14336_ clknet_leaf_56_clk _01449_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfxtp_1
Xhold508 cpu.RF0.registers\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold519 cpu.RF0.registers\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ clknet_leaf_13_clk _01380_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ net1760 net201 net375 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09377__A0 _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ clknet_leaf_95_clk _00398_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09328__A _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ clknet_leaf_59_clk _01311_ net1348 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10526__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13149_ clknet_leaf_52_clk _00329_ net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1208 cpu.RF0.registers\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 cpu.RF0.registers\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_07710_ net1033 cpu.RF0.registers\[18\]\[17\] net769 vssd1 vssd1 vccd1 vccd1 _03001_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13628__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ cpu.RF0.registers\[8\]\[1\] _02014_ net685 cpu.RF0.registers\[24\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07641_ cpu.RF0.registers\[24\]\[13\] net608 _02906_ _02913_ _02922_ vssd1 vssd1
+ vccd1 vccd1 _02932_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09998__A cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07572_ _02851_ _02854_ _02855_ _02856_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ _03407_ _04205_ _04553_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__and3_1
X_06523_ cpu.f0.num\[19\] net1020 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__xor2_1
XANTENNA__10998__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _04430_ _04439_ net450 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ net2858 _01841_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__nor2_1
XANTENNA__07863__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13008__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12574__D cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ net468 _03931_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__nor2_1
X_06385_ cpu.f0.num\[11\] vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08407__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ net1078 cpu.RF0.registers\[30\]\[23\] net837 vssd1 vssd1 vccd1 vccd1 _03415_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06969__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ net943 cpu.RF0.registers\[11\]\[25\] net879 vssd1 vssd1 vccd1 vccd1 _03346_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ net1028 cpu.RF0.registers\[19\]\[23\] net820 vssd1 vssd1 vccd1 vccd1 _02297_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13158__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout593_A _02162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14403__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08040__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1300_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ cpu.RF0.registers\[11\]\[26\] net690 net674 cpu.RF0.registers\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout760_A _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09244__Y _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ cpu.RF0.registers\[0\]\[30\] net617 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14553__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ cpu.RF0.registers\[11\]\[17\] net690 _04166_ _04173_ _04175_ vssd1 vssd1
+ vccd1 vccd1 _04179_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_51_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ cpu.RF0.registers\[24\]\[24\] net607 net566 cpu.RF0.registers\[11\]\[24\]
+ _03129_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a221o_1
XANTENNA__08894__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__B2 cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ net2163 net228 net431 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06884__X _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09509_ _04798_ _04799_ net486 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10781_ net287 _05732_ _05733_ net1016 cpu.IM0.address_IM\[19\] vssd1 vssd1 vccd1
+ vccd1 _05734_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12520_ _06294_ _06295_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08317__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__Q cpu.IM0.address_IM\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12451_ _01887_ _01942_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11402_ net2056 net236 net385 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12382_ net1119 net1654 net529 net1036 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ clknet_leaf_105_clk _01234_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11333_ net2795 net138 net394 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
XANTENNA__12126__X _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ clknet_leaf_97_clk _01165_ net1231 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14083__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ net2274 net147 net404 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__mux2_1
XANTENNA__08052__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07594__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ clknet_leaf_43_clk _00192_ net1303 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
X_10215_ cpu.IM0.address_IM\[31\] net930 _05475_ _05476_ vssd1 vssd1 vccd1 vccd1 _00054_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08031__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ net2717 net159 net411 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__mux2_1
XANTENNA__08987__A _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ net125 _05413_ _05410_ net625 vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11617__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__Y _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09531__A0 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07137__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ clknet_leaf_77_clk _01018_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13920__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ clknet_leaf_74_clk _00949_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14069__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08098__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ clknet_leaf_78_clk _00880_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ net282 _05870_ net986 vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11352__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__B2 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12718_ net1475 cpu.LCD0.row_2\[112\] net1010 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__mux2_1
XANTENNA__07845__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10476__B net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13698_ clknet_leaf_95_clk _00811_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07769__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10995__A3 _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ net2551 net2512 net999 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12197__A2 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10974__A_N _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold305 cpu.RF0.registers\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ clknet_leaf_57_clk _01432_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold316 cpu.RF0.registers\[24\]\[4\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 cpu.FetchedInstr\[8\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 cpu.RF0.registers\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 cpu.LCD0.row_2\[75\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09860_ cpu.IM0.address_IM\[2\] _02644_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__xnor2_1
Xfanout807 net808 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_2
XANTENNA__13450__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14576__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net819 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
Xfanout829 _02129_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
X_08811_ net1083 cpu.RF0.registers\[16\]\[19\] net841 vssd1 vssd1 vccd1 vccd1 _04102_
+ sky130_fd_sc_hd__and3_1
X_09791_ _04605_ _04885_ net478 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__mux2_1
Xhold1005 cpu.RF0.registers\[18\]\[4\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11527__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1016 cpu.RF0.registers\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03902_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nand2b_1
Xhold1027 cpu.LCD0.row_1\[58\] vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 cpu.RF0.registers\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12212__A _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1049 cpu.LCD0.row_2\[42\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_clk_X clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ cpu.IM0.address_IM\[2\] net554 _03962_ _03963_ vssd1 vssd1 vccd1 vccd1 _03964_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_75_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07624_ net964 cpu.RF0.registers\[10\]\[13\] net786 vssd1 vssd1 vccd1 vccd1 _02915_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07025__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__A_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ net970 cpu.RF0.registers\[2\]\[8\] net771 vssd1 vssd1 vccd1 vccd1 _02846_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout341_A _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__Y _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__B net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ cpu.f0.num\[16\] cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07836__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ net1060 cpu.RF0.registers\[22\]\[5\] net802 vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07679__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07300__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ net511 _04294_ _04453_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__o31a_1
X_06437_ _01844_ _01845_ net2851 vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[16\] sky130_fd_sc_hd__mux2_1
XFILLER_0_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10954__X _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1250_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_A _02144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_12_clk_X clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ net511 _04363_ _04364_ _04445_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__o31ai_4
X_06368_ cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06880__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08107_ cpu.RF0.registers\[23\]\[22\] net671 net651 cpu.RF0.registers\[7\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__a22o_1
XANTENNA__10606__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ _02113_ _02117_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__nor2_1
XANTENNA__08261__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ cpu.RF0.registers\[20\]\[24\] net709 net658 cpu.RF0.registers\[13\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold850 cpu.RF0.registers\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _01701_ vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_X clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold872 cpu.DM0.readdata\[6\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _00241_ vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold894 cpu.RF0.registers\[21\]\[14\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ cpu.IM0.address_IM\[12\] _02869_ _02904_ cpu.IM0.address_IM\[13\] vssd1 vssd1
+ vccd1 vccd1 _05279_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09989_ _05267_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13943__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A2 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12112__A2 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ net1788 net169 net319 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__mux2_1
XANTENNA__08867__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ net738 _05131_ _05820_ _02001_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a211o_1
X_14670_ net1392 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
X_11882_ net1950 net187 net328 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ cpu.IM0.address_IM\[1\] _05771_ net721 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__mux2_4
X_13621_ clknet_leaf_73_clk _00734_ net1341 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06774__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ net2755 net561 net536 _05721_ vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__a22o_1
X_13552_ clknet_leaf_75_clk _00665_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07589__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10296__B cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13323__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14449__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ _01811_ _06284_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13483_ clknet_leaf_89_clk _00596_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ cpu.LCD0.row_1\[101\] cpu.LCD0.row_1\[109\] net899 vssd1 vssd1 vccd1 vccd1
+ _00325_ sky130_fd_sc_hd__mux2_1
XANTENNA__12179__A2 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ cpu.DM0.data_i\[25\] net534 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__and2_1
XANTENNA__10583__Y _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ net1123 net2677 net531 cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 _01491_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_101_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13473__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ clknet_leaf_7_clk _01217_ net1162 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11316_ net2257 net198 net395 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ cpu.LCD0.row_1\[127\] _06014_ _06179_ _06189_ net556 vssd1 vssd1 vccd1 vccd1
+ _06190_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_82_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ clknet_leaf_68_clk _01148_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11247_ net1741 net202 net403 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__mux2_1
XANTENNA__08004__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net2646 net223 net413 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__mux2_1
XANTENNA__08510__A _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10129_ _05395_ _05397_ _05392_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_66_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09504__A0 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09044__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_92_clk _00932_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09807__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06684__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ cpu.RF0.registers\[21\]\[3\] net593 _02608_ _02614_ _02617_ vssd1 vssd1 vccd1
+ vccd1 _02631_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07271_ net980 cpu.RF0.registers\[7\]\[7\] net818 vssd1 vssd1 vccd1 vccd1 _02562_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_73_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08491__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09010_ net934 cpu.RF0.registers\[1\]\[31\] net882 vssd1 vssd1 vccd1 vccd1 _04301_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11810__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 cpu.f0.data_adr\[27\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _00161_ vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _01718_ vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 net75 vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A2 _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 cpu.SR1.char_in\[3\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 cpu.RF0.registers\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13966__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold168 cpu.RF0.registers\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ cpu.IM0.address_IM\[6\] _05189_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__xor2_1
Xhold179 _01625_ vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10950__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 _02146_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_6
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_6
Xfanout626 _02101_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09743__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _04573_ _04872_ net480 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__mux2_1
Xfanout637 _02066_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_84_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10353__A1 _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 _02059_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_8
XANTENNA__08420__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12213__Y _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__B2 cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _02054_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11257__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12990__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _04399_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__and2_1
X_06986_ net1028 cpu.RF0.registers\[18\]\[23\] net769 vssd1 vssd1 vccd1 vccd1 _02277_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07036__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ cpu.RF0.registers\[31\]\[0\] net1096 net857 vssd1 vssd1 vccd1 vccd1 _04016_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08849__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1298_A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08656_ net1102 cpu.RF0.registers\[17\]\[2\] net884 vssd1 vssd1 vccd1 vccd1 _03947_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09889__C cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07607_ net1046 cpu.RF0.registers\[30\]\[12\] net764 net831 cpu.RF0.registers\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ net1101 cpu.RF0.registers\[20\]\[4\] net876 vssd1 vssd1 vccd1 vccd1 _03878_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout723_A _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _02825_ _02827_ _02828_ _02798_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o31a_4
XTAP_TAPCELL_ROW_46_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09274__A2 _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07469_ net482 net471 net468 _02756_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__Y _02172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ net441 net439 net461 vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__mux2_1
X_10480_ net1516 net922 net747 a1.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__a22o_1
XANTENNA__09026__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__B _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10263__C_N net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _04428_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08234__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12150_ cpu.LCD0.row_2\[121\] _06022_ _06024_ cpu.LCD0.row_1\[97\] vssd1 vssd1 vccd1
+ vccd1 _06050_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ cpu.RF0.registers\[2\]\[31\] net128 net422 vssd1 vssd1 vccd1 vccd1 _00535_
+ sky130_fd_sc_hd__mux2_1
X_12081_ cpu.LCD0.nextState\[3\] cpu.LCD0.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _05982_
+ sky130_fd_sc_hd__nor2_4
Xhold680 cpu.RF0.registers\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 cpu.f0.num\[28\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08968__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _05906_ _05907_ cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11167__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ clknet_leaf_44_clk net1506 net1305 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10859__X _05790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1380 cpu.RF0.registers\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1391 cpu.RF0.registers\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
X_11934_ net2215 net241 net320 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14271__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ clknet_leaf_54_clk _01754_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11865_ net2807 net255 net329 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
X_13604_ clknet_leaf_99_clk _00717_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ net1612 net560 net538 _05758_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14584_ clknet_leaf_53_clk net2200 net1363 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_11796_ net2772 net131 net338 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ clknet_leaf_105_clk _00648_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10747_ net992 _04830_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11630__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10280__B1 cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ cpu.LCD0.row_1\[84\] cpu.LCD0.row_1\[92\] net903 vssd1 vssd1 vccd1 vccd1
+ _00308_ sky130_fd_sc_hd__mux2_1
XANTENNA__09017__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13466_ clknet_leaf_97_clk _00579_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10754__B _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13989__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net1548 net730 net501 _06232_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__o22a_1
X_13397_ clknet_leaf_73_clk _00510_ net1341 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12348_ cpu.LCD0.cnt_20ms\[15\] cpu.LCD0.cnt_20ms\[14\] _06212_ cpu.LCD0.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06787__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12279_ cpu.LCD0.row_1\[15\] _05994_ _06001_ cpu.LCD0.row_1\[71\] _06172_ vssd1 vssd1
+ vccd1 vccd1 _06173_ sky130_fd_sc_hd__a221o_1
X_14018_ clknet_leaf_95_clk _01131_ net1219 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08878__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06840_ net1067 net1065 net1072 net1069 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_88_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13369__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06771_ net1111 net1113 net1114 net1117 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__and4bb_4
XANTENNA__14614__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08510_ _03797_ _03800_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nor2_1
XANTENNA__11805__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ _04760_ _04780_ net456 vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__mux2_1
XANTENNA__07503__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08700__A1 cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _03729_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nand2_1
XANTENNA__09071__A _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08372_ cpu.RF0.registers\[0\]\[11\] net662 net548 vssd1 vssd1 vccd1 vccd1 _03663_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload76_A clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08118__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ net975 cpu.RF0.registers\[15\]\[3\] net829 vssd1 vssd1 vccd1 vccd1 _02614_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11540__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07254_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__inv_2
XANTENNA__10810__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07957__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__Q a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06861__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07019__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__B1 _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ net969 cpu.RF0.registers\[5\]\[10\] net797 vssd1 vssd1 vccd1 vccd1 _02476_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1046_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10574__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14144__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout401 _05921_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_8
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _03436_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout673_A _02042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 net459 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ net511 _04665_ _05108_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__o31ai_4
Xfanout467 net469 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
Xfanout478 net483 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07742__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14294__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net459 _05019_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout840_A _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06969_ cpu.RF0.registers\[5\]\[25\] net603 net576 cpu.RF0.registers\[14\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout938_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ cpu.RF0.registers\[11\]\[0\] net688 net681 cpu.RF0.registers\[18\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _04710_ _04972_ _04977_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_48_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ cpu.RF0.registers\[0\]\[3\] net663 net550 vssd1 vssd1 vccd1 vccd1 _03930_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14684__1406 vssd1 vssd1 vccd1 vccd1 _14684__1406/HI net1406 sky130_fd_sc_hd__conb_1
X_11650_ net1621 net189 net354 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XANTENNA__12886__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11015__B1_N net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ cpu.LCD0.row_1\[7\] net2178 net904 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XANTENNA__08028__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ net2293 net196 net364 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__mux2_1
XANTENNA__08455__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11450__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ net1132 net2331 net912 _05653_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_94_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13320_ clknet_leaf_21_clk cpu.RU0.next_FetchedData\[27\] net1173 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06481__A2 _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13251_ clknet_leaf_27_clk _00431_ net1188 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08207__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ net12 net754 net564 a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12202_ _06093_ _06095_ _06097_ _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ clknet_leaf_36_clk _00362_ net1265 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07415__D1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10394_ cpu.f0.i\[9\] net271 vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
X_12133_ _05981_ _05995_ _05997_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__and3_4
X_12064_ cpu.LCD0.cnt_500hz\[9\] _05969_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__and2_1
XANTENNA__10317__A1 cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13511__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14637__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _02207_ net532 net282 vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__o21ba_1
Xfanout990 net996 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09443__X _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__X _05683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13661__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ clknet_leaf_44_clk net1514 net1306 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ net2919 net182 net323 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08694__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12897_ clknet_leaf_27_clk _00086_ net1189 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ clknet_leaf_26_clk _01737_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11848_ net1772 net190 net330 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XANTENNA__14017__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08446__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ clknet_leaf_56_clk _01669_ net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_11779_ net2485 net193 net340 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__mux2_1
XANTENNA__11360__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13518_ clknet_leaf_5_clk _00631_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14498_ clknet_leaf_51_clk _01600_ net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload11 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_2
X_13449_ clknet_leaf_104_clk _00562_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload22 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14167__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload33 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_6
Xclkload44 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload44/X sky130_fd_sc_hd__clkbuf_4
Xclkload55 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_16
XANTENNA__09946__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload66 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10556__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload77 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_8
Xclkload88 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload99 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__inv_6
X_08990_ _03371_ _03373_ _03337_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a21o_1
XANTENNA__13191__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07972__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ cpu.CU0.bit30 net633 net519 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a21o_1
X_07872_ cpu.RF0.registers\[10\]\[28\] net570 _03162_ net623 vssd1 vssd1 vccd1 vccd1
+ _03163_ sky130_fd_sc_hd__a211o_1
XANTENNA__10005__A cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net468 _04898_ _04901_ net290 _04900_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o221a_1
X_06823_ net1118 _02082_ _02083_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__and3_1
XANTENNA__11535__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09513__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ _04421_ _04424_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__nor2_1
X_06754_ net1096 net845 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06856__C net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ net482 _04758_ _04763_ _04695_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__o211a_1
XANTENNA__08685__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ net1825 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[21\] sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_90_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10492__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ cpu.RF0.registers\[27\]\[9\] net711 net702 cpu.RF0.registers\[5\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08355_ net941 cpu.RF0.registers\[7\]\[11\] net847 vssd1 vssd1 vccd1 vccd1 _03646_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08437__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ cpu.RF0.registers\[5\]\[4\] net602 net590 cpu.RF0.registers\[15\]\[4\] _02596_
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_A _02210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_74_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08286_ net1086 cpu.RF0.registers\[19\]\[13\] net835 vssd1 vssd1 vccd1 vccd1 _03577_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10394__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__A1 cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07237_ net955 cpu.RF0.registers\[5\]\[9\] net795 vssd1 vssd1 vccd1 vccd1 _02528_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1330_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07984__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ cpu.RF0.registers\[16\]\[11\] net582 _02449_ _02451_ _02456_ vssd1 vssd1
+ vccd1 vccd1 _02459_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout790_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07099_ net1049 cpu.RF0.registers\[21\]\[14\] net797 vssd1 vssd1 vccd1 vccd1 _02390_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07963__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1209 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_4
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net223 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout1229 net1232 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout231 _05783_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net244 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08311__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 net267 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13684__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08912__A1 _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 _04393_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ net478 _04744_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__nor2_1
XANTENNA__11445__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ clknet_leaf_15_clk _00039_ net1243 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09423__B _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07224__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__Q cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12751_ net1498 net496 net281 cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_81_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08140__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10483__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11702_ net1985 net247 net347 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12682_ cpu.LCD0.row_2\[84\] cpu.LCD0.row_2\[76\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ clknet_leaf_17_clk _01532_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11027__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11633_ net1678 net238 net357 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
XANTENNA__08428__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13064__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12129__X _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11180__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14352_ clknet_leaf_57_clk _01465_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11564_ net2917 net138 net366 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
XANTENNA__07597__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13303_ clknet_leaf_31_clk cpu.RU0.next_FetchedData\[10\] net1206 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[10\] sky130_fd_sc_hd__dfrtp_1
X_10515_ net62 net918 vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__and2_1
X_11495_ net1644 net150 net375 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
X_14283_ clknet_leaf_90_clk _01396_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10446_ net24 net754 net564 a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__a22o_1
X_13234_ clknet_leaf_44_clk _00414_ net1304 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10538__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__Y _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13165_ clknet_leaf_37_clk _00345_ net1263 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_10377_ net1126 _05606_ net266 net2074 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08600__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12901__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12116_ cpu.LCD0.row_1\[0\] _06015_ _06016_ cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1
+ vccd1 _06017_ sky130_fd_sc_hd__a22o_1
X_13096_ clknet_leaf_49_clk _00276_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09156__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _01954_ _05957_ _05960_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__and3_1
XANTENNA__07118__B _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A1 cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11355__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ clknet_leaf_1_clk _01111_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13658__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08667__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09052__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ clknet_leaf_20_clk _00138_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13407__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10474__B1 _05640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08131__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06470_ cpu.DM0.state\[1\] cpu.DM0.state\[2\] cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1
+ _01866_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14619_ clknet_leaf_29_clk _01720_ net1203 vssd1 vssd1 vccd1 vccd1 cpu.RU0.InstrRead
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11018__A2 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09616__C1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06692__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11090__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08140_ cpu.RF0.registers\[27\]\[23\] net711 net670 cpu.RF0.registers\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a22o_1
XANTENNA__10777__A1 cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13557__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08071_ cpu.RF0.registers\[18\]\[25\] net680 _03341_ _03342_ _03343_ vssd1 vssd1
+ vccd1 vccd1 _03362_ sky130_fd_sc_hd__a2111o_1
Xclkload100 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07022_ net742 net741 _02091_ net628 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1
+ _02313_ sky130_fd_sc_hd__o41a_4
XANTENNA_wire856_A _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload39_A clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14683__1405 vssd1 vssd1 vccd1 vccd1 _14683__1405/HI net1405 sky130_fd_sc_hd__conb_1
X_08973_ cpu.RF0.registers\[10\]\[26\] net691 _04249_ _04256_ _04258_ vssd1 vssd1
+ vccd1 vccd1 _04264_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 cpu.LCD0.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 cpu.FetchedInstr\[5\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ net957 cpu.RF0.registers\[11\]\[30\] net776 vssd1 vssd1 vccd1 vccd1 _03215_
+ sky130_fd_sc_hd__and3_1
Xhold39 cpu.f0.write_data\[10\] vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07855_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08370__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06806_ _02096_ _01778_ _02091_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07786_ _03073_ _03075_ _03076_ _03046_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__o31a_1
XFILLER_0_79_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _02507_ _03698_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__nand2_1
X_06737_ net943 net879 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__and2_2
XANTENNA__13087__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10465__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ a1.CPU_DAT_O\[4\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[4\]
+ sky130_fd_sc_hd__and2_1
X_09456_ net298 _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09870__A2 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11009__A2 _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ cpu.IM0.address_IM\[10\] net554 _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__a22o_4
X_09387_ net472 _04440_ _04567_ _04673_ _04676_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ _01757_ _01968_ _01758_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1166_X net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08338_ cpu.IM0.address_IM\[12\] net552 _03627_ _03628_ vssd1 vssd1 vccd1 vccd1 _03629_
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10768__A1 a1.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08269_ cpu.RF0.registers\[31\]\[15\] net686 net657 cpu.RF0.registers\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a22o_1
XANTENNA__12924__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ net527 _05538_ _05542_ _05541_ net728 vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a311o_2
XFILLER_0_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net2107 net212 net399 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _01798_ net307 _05482_ _05483_ net728 vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a221o_2
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07936__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ cpu.IM0.address_IM\[27\] _02211_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1004 net1012 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_2
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10940__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 net1033 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_2
XFILLER_0_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10093_ cpu.IM0.address_IM\[21\] _05355_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__xnor2_2
Xfanout1037 cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_2
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1059 net1064 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07506__X _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09434__A _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ clknet_leaf_63_clk _01034_ net1309 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11175__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ clknet_leaf_8_clk _00965_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12803_ net2255 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10867__X _05796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13783_ clknet_leaf_64_clk _00896_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10995_ net274 _05881_ _05882_ net926 net2857 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__a32o_1
XANTENNA__09846__C1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11903__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _06316_ _01762_ _01764_ net498 cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1
+ _01721_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__Y _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12665_ net2399 net2338 net998 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__mux2_1
XANTENNA__10208__B1 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14404_ clknet_leaf_23_clk _01515_ net1194 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_11616_ net1685 net206 net358 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09074__A0 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12596_ _01757_ _01755_ _01985_ _01758_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a31o_1
X_14335_ clknet_leaf_51_clk _01448_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08821__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ net1640 net197 net366 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07828__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 cpu.RF0.registers\[4\]\[3\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ clknet_leaf_93_clk _01379_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08513__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ net1984 net212 net375 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XANTENNA__09377__A1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ clknet_leaf_99_clk _00397_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ net1124 _05632_ net265 net2261 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__a2bb2o_1
X_14197_ clknet_leaf_74_clk _01310_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07388__B1 _02676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07927__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ clknet_leaf_50_clk _00328_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09047__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14205__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ clknet_leaf_46_clk net2390 net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1209 cpu.RF0.registers\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11085__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ cpu.RF0.registers\[13\]\[13\] net597 _02905_ _02907_ _02910_ vssd1 vssd1
+ vccd1 vccd1 _02931_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14355__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07560__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ cpu.RF0.registers\[8\]\[8\] net612 _02848_ net623 vssd1 vssd1 vccd1 vccd1
+ _02862_ sky130_fd_sc_hd__a211o_1
XANTENNA__09998__B _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08104__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06522_ cpu.f0.num\[0\] cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__xor2_1
XANTENNA__11813__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ net512 _04579_ _04580_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o31a_2
XFILLER_0_53_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10998__A1 a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06453_ _01841_ _01856_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[11\] sky130_fd_sc_hd__nor2_1
XFILLER_0_29_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _04530_ _04531_ net476 vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12947__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _04456_ _04462_ net473 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__mux2_1
X_06384_ cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09604__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ net1078 cpu.RF0.registers\[25\]\[23\] net862 vssd1 vssd1 vccd1 vccd1 _03414_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08126__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07030__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11401__X _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ net1087 cpu.RF0.registers\[19\]\[25\] _02062_ vssd1 vssd1 vccd1 vccd1 _03345_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_86_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14280__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12941__Q a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ net955 cpu.RF0.registers\[1\]\[23\] net804 vssd1 vssd1 vccd1 vccd1 _02296_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09368__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09368__B2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07039__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08956_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__inv_2
XANTENNA__06878__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07907_ net488 _03195_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__o21ai_1
X_08887_ cpu.RF0.registers\[29\]\[17\] net672 net671 cpu.RF0.registers\[23\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ cpu.RF0.registers\[23\]\[24\] net614 net602 cpu.RF0.registers\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
XANTENNA__13722__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ net1039 cpu.RF0.registers\[20\]\[21\] net781 vssd1 vssd1 vccd1 vccd1 _03060_
+ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_36_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1283_X net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09508_ _04738_ _04740_ net476 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__mux2_1
XANTENNA__09701__B _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10780_ net986 cpu.f0.data_adr\[19\] vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__or2_2
XFILLER_0_71_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10989__A1 _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07303__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09439_ _04566_ _04654_ _04658_ net272 _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07854__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ cpu.DM0.dhit cpu.f0.i\[0\] _06249_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _05766_ _05906_ net503 vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__and3_4
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12554__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ net1119 net2330 net529 net1065 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14120_ clknet_leaf_98_clk _01233_ net1232 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11332_ net2629 net143 net397 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
XANTENNA__13102__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07082__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14228__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ clknet_leaf_77_clk _01164_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ net1906 net150 net403 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13002_ clknet_leaf_43_clk _00191_ net1303 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
X_10214_ net628 _04446_ net931 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a21oi_1
X_11194_ net1937 net180 net412 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__mux2_1
XANTENNA__13252__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08582__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _05411_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__nor2_1
XANTENNA__14378__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _05325_ _05336_ _05335_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a21o_1
XANTENNA__09531__A1 _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08334__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13904_ clknet_leaf_73_clk _01017_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13835_ clknet_leaf_91_clk _00948_ net1278 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_27_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11633__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ clknet_leaf_6_clk _00879_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09295__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10978_ _02981_ net532 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12717_ cpu.LCD0.row_2\[119\] net2439 net1006 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__mux2_1
XANTENNA__07845__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682__1404 vssd1 vssd1 vccd1 vccd1 _14682__1404/HI net1404 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_80_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13697_ clknet_leaf_67_clk _00810_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12648_ net2502 net2455 net999 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09598__A1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12579_ _06325_ _06337_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__and2b_2
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10601__A0 cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14318_ clknet_leaf_0_clk _01431_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold306 a1.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 cpu.RF0.registers\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold328 cpu.RF0.registers\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 a1.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ clknet_leaf_106_clk _01362_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10365__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout819 _02134_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
X_08810_ net1085 cpu.RF0.registers\[23\]\[19\] net844 vssd1 vssd1 vccd1 vccd1 _04101_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11808__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _02410_ _03535_ _05080_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__a21oi_1
Xhold1006 cpu.LCD0.row_2\[24\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 cpu.RF0.registers\[18\]\[18\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _03899_ _03901_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__or2_1
Xhold1028 cpu.RF0.registers\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 cpu.RF0.registers\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08325__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ cpu.RF0.registers\[0\]\[2\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03963_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07623_ net1045 cpu.RF0.registers\[25\]\[13\] net757 vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11543__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout167_A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13895__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__B _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__X _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ net1052 cpu.RF0.registers\[25\]\[8\] net759 vssd1 vssd1 vccd1 vccd1 _02845_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09286__B1 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08418__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07322__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06505_ cpu.f0.num\[27\] cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07485_ net982 cpu.RF0.registers\[5\]\[5\] net798 vssd1 vssd1 vccd1 vccd1 _02776_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout334_A _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ _04514_ _04494_ _04490_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__and3b_2
XFILLER_0_91_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06436_ net1908 _01842_ _01845_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[15\] sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13125__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09589__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06367_ net1095 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__inv_2
X_09155_ net511 _04363_ _04364_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1243_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06880__B net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08106_ _03393_ _03394_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_40_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07695__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ net449 _04373_ _04375_ _04376_ net301 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13275__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08037_ _03324_ _03325_ _03326_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 cpu.RF0.registers\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14520__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1129_X net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 cpu.RF0.registers\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07992__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 cpu.RF0.registers\[27\]\[9\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 cpu.RF0.registers\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09210__A0 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold884 cpu.RF0.registers\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 cpu.RF0.registers\[15\]\[14\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11718__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10622__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ cpu.IM0.address_IM\[12\] _02869_ _05259_ _05261_ vssd1 vssd1 vccd1 vccd1
+ _05268_ sky130_fd_sc_hd__a22o_1
XANTENNA__07056__X _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ cpu.RF0.registers\[4\]\[27\] net677 _04216_ _04226_ _04227_ vssd1 vssd1 vccd1
+ vccd1 _04230_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06401__A cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ net2777 net181 net321 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06895__X _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11320__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09712__A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ cpu.DM0.readdata\[21\] net734 vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ net2218 net189 net326 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11453__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ clknet_leaf_71_clk _00733_ net1340 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ cpu.DM0.readdata\[1\] _05058_ net739 vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12846__Q cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07232__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07827__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ clknet_leaf_82_clk _00664_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10763_ cpu.IM0.address_IM\[14\] net1017 net284 _05720_ vssd1 vssd1 vccd1 vccd1 _05721_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ net262 _06283_ _06284_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13482_ clknet_leaf_100_clk _00595_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ cpu.LCD0.row_1\[100\] cpu.LCD0.row_1\[108\] net903 vssd1 vssd1 vccd1 vccd1
+ _00324_ sky130_fd_sc_hd__mux2_1
X_12433_ cpu.DM0.readdata\[24\] net730 net500 _06240_ vssd1 vssd1 vccd1 vccd1 _01540_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ net1122 net1770 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08063__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14103_ clknet_leaf_65_clk _01216_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11315_ net2689 net211 net395 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__mux2_1
X_12295_ _06181_ _06183_ _06185_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__or4_1
X_14034_ clknet_leaf_59_clk _01147_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ net2397 net213 net402 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__mux2_1
XANTENNA__13768__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11628__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10898__A0 cpu.DM0.readdata\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ net2191 net224 net412 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__mux2_1
X_10128_ _05369_ _05381_ _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09504__A1 _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ net626 _05117_ net1023 vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_86_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ clknet_leaf_92_clk _00931_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09268__B1 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13148__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13749_ clknet_leaf_73_clk _00862_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07270_ net980 cpu.RF0.registers\[3\]\[7\] net823 vssd1 vssd1 vccd1 vccd1 _02561_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07294__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13298__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09069__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07046__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__A1 cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold103 net91 vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold114 net79 vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 cpu.f0.write_data\[27\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _00163_ vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold147 cpu.RF0.registers\[0\]\[19\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 cpu.RF0.registers\[27\]\[11\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _05195_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__xnor2_1
Xhold169 cpu.RF0.registers\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10338__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10950__B _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload21_A clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout605 _02144_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_6
XANTENNA__09743__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _02132_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11538__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _03568_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__xnor2_2
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_2
Xfanout638 _02065_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_6
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06557__A1 cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout649 _02058_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_52_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07317__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _04543_ _04758_ net479 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__mux2_1
X_06985_ net1028 cpu.RF0.registers\[25\]\[23\] net756 vssd1 vssd1 vccd1 vccd1 _02276_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout284_A _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ cpu.RF0.registers\[25\]\[0\] net1096 net863 vssd1 vssd1 vccd1 vccd1 _04015_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10949__Y _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ cpu.RF0.registers\[12\]\[2\] net697 _03943_ _03944_ _03945_ vssd1 vssd1 vccd1
+ vccd1 _03946_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout451_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11273__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ cpu.RF0.registers\[15\]\[12\] net590 _02875_ _02877_ _02887_ vssd1 vssd1
+ vccd1 vccd1 _02897_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08586_ net1100 cpu.RF0.registers\[19\]\[4\] net836 vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_77_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ _02816_ _02818_ _02819_ _02820_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07987__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07285__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ net481 net472 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ net300 _04158_ net469 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__mux2_1
X_06419_ cpu.c0.count\[8\] cpu.c0.count\[11\] cpu.c0.count\[9\] vssd1 vssd1 vccd1
+ vccd1 _01832_ sky130_fd_sc_hd__or3b_1
XFILLER_0_84_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07399_ cpu.RF0.registers\[11\]\[0\] net566 _02687_ _02688_ _02689_ vssd1 vssd1 vccd1
+ vccd1 _02690_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09138_ net467 _03899_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08314__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13910__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ net438 _04358_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10592__A2 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ net2850 net137 net422 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__mux2_1
XANTENNA__07993__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ cpu.LCD0.nextState\[0\] cpu.LCD0.nextState\[1\] vssd1 vssd1 vccd1 vccd1 _05981_
+ sky130_fd_sc_hd__and2b_2
XANTENNA__08611__A _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 cpu.RF0.registers\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 cpu.RF0.registers\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08537__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 cpu.RF0.registers\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11448__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ cpu.IG0.Instr\[10\] cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nor2_2
X_14681__1403 vssd1 vssd1 vccd1 vccd1 _14681__1403/HI net1403 sky130_fd_sc_hd__conb_1
XANTENNA__06769__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_36_clk _00171_ net1303 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1370 cpu.RF0.registers\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1381 cpu.LCD0.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14416__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ net1974 net245 net320 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
Xhold1392 cpu.DM0.readdata\[4\] vssd1 vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11183__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ clknet_leaf_54_clk _01753_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11864_ net1836 net239 net329 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
X_13603_ clknet_leaf_78_clk _00716_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10815_ cpu.IM0.address_IM\[29\] net1014 net285 _05757_ vssd1 vssd1 vccd1 vccd1 _05758_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14583_ clknet_leaf_56_clk net2453 net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_11795_ net1713 net136 net338 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14566__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13440__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ clknet_leaf_85_clk _00647_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10746_ net2409 net560 net538 _05708_ vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13465_ clknet_leaf_42_clk _00578_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10677_ net1819 cpu.LCD0.row_1\[91\] net898 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
X_12416_ cpu.DM0.data_i\[16\] net535 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_73_clk_X clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13396_ clknet_leaf_72_clk _00509_ net1340 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13590__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12347_ net1507 _06213_ _06215_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08080__X _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12278_ cpu.LCD0.row_2\[103\] _06018_ _06031_ cpu.LCD0.row_1\[31\] vssd1 vssd1 vccd1
+ vccd1 _06172_ sky130_fd_sc_hd__a22o_1
XANTENNA__08521__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11358__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__A2 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ clknet_leaf_64_clk _01130_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11229_ net1996 net155 net406 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_clk_X clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06539__B2 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09055__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06770_ net1092 net865 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_11_clk_X clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14096__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11093__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08440_ _02544_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_clk_X clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08371_ _03651_ _03653_ _03658_ _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07322_ net1063 cpu.RF0.registers\[20\]\[3\] net782 vssd1 vssd1 vccd1 vccd1 _02613_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__B1 _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A2 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13933__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload69_A clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07253_ net546 _02543_ _02509_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a21o_2
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08216__A1 _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ cpu.RF0.registers\[0\]\[10\] net619 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__or2_1
XANTENNA__07019__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__A1 cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1039_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout499_A _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _05919_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout413 _05917_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1206_A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
Xfanout446 _03335_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _05115_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__inv_2
Xfanout457 net459 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13313__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14439__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_2
Xfanout479 net483 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_2
XANTENNA_fanout666_A _02050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09756_ net459 _04874_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__or2_1
XANTENNA__10900__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ cpu.RF0.registers\[8\]\[25\] net611 net593 cpu.RF0.registers\[21\]\[25\]
+ _02251_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a221o_1
XANTENNA__06886__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ cpu.RF0.registers\[27\]\[0\] net712 net692 cpu.RF0.registers\[10\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__a22o_1
X_09687_ net471 _03964_ _04974_ _03931_ net482 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__o32ai_1
XTAP_TAPCELL_ROW_48_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ net966 net787 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__and2_1
XANTENNA__08152__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14589__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _03918_ _03920_ _03925_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__or4_1
XANTENNA__10201__A cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ cpu.RF0.registers\[17\]\[5\] net694 net669 cpu.RF0.registers\[22\]\[5\] _03842_
+ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1363_X net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10600_ cpu.LCD0.row_1\[6\] net2336 net908 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ net2070 net197 net362 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12251__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10531_ net41 net918 vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_94_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06856__A_N net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ clknet_leaf_23_clk _00430_ net1177 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09404__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ net11 net754 net564 net2816 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ cpu.LCD0.row_1\[83\] _05986_ _06018_ cpu.LCD0.row_2\[99\] _06098_ vssd1 vssd1
+ vccd1 vccd1 _06099_ sky130_fd_sc_hd__a221o_1
X_13181_ clknet_leaf_30_clk _00361_ net1207 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10393_ net1125 _05614_ net267 net2128 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12132_ net746 _05982_ _05996_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__and3_4
XANTENNA__11178__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ cpu.LCD0.cnt_500hz\[9\] _05969_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__or2_1
XANTENNA__11514__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net1918 net925 net273 _05895_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08391__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
Xfanout991 net994 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07733__A3 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13806__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ clknet_leaf_44_clk net1465 net1305 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14663__1387 vssd1 vssd1 vccd1 vccd1 _14663__1387/HI net1387 sky130_fd_sc_hd__conb_1
X_11916_ net1776 _05817_ net322 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07497__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10111__A cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ clknet_leaf_28_clk _00010_ net1188 vssd1 vssd1 vccd1 vccd1 a1.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14635_ clknet_leaf_31_clk _01736_ net1206 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13956__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ net2066 net206 net330 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
XANTENNA__12737__S _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11641__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14566_ clknet_leaf_47_clk _01668_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[77\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07249__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__A2 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ net1774 net199 net339 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__mux2_1
XANTENNA__10765__B _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08516__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ clknet_leaf_101_clk _00630_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ net2842 net559 net537 _05696_ vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14497_ clknet_leaf_49_clk _01599_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12980__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13448_ clknet_leaf_98_clk _00561_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_49_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload34 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_8
Xclkload45 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload45/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09946__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload56 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_16
X_13379_ clknet_leaf_77_clk _00492_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload67 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinv_4
Xclkload78 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_80_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11753__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload89 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_clkbuf_leaf_53_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13336__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11088__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ cpu.CU0.bit30 net633 net519 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a21oi_1
X_07871_ net1050 cpu.RF0.registers\[31\]\[28\] net830 net581 cpu.RF0.registers\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a32o_1
X_09610_ net463 _04025_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__nor2_1
XANTENNA__11816__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ cpu.CU0.funct3\[0\] _02107_ _02083_ _01846_ vssd1 vssd1 vccd1 vccd1 _02113_
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__13486__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _03735_ _03769_ _04040_ net513 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06753_ net1110 net1112 net1114 net1116 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__and4b_1
X_09472_ net487 _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__or2_1
XANTENNA__06856__D net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__A cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06684_ net1422 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[20\] sky130_fd_sc_hd__and2_1
XANTENNA__12481__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ net935 cpu.RF0.registers\[12\]\[9\] net867 vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07033__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _05776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ net1087 cpu.RF0.registers\[22\]\[11\] net851 vssd1 vssd1 vccd1 vccd1 _03645_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06872__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14680__1402 vssd1 vssd1 vccd1 vccd1 _14680__1402/HI net1402 sky130_fd_sc_hd__conb_1
X_07305_ cpu.RF0.registers\[27\]\[4\] net592 net575 cpu.RF0.registers\[14\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XANTENNA__07330__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12944__Q a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload6 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinv_4
X_08285_ net1086 cpu.RF0.registers\[27\]\[13\] net880 vssd1 vssd1 vccd1 vccd1 _03576_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout414_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ net1034 cpu.RF0.registers\[22\]\[9\] net799 vssd1 vssd1 vccd1 vccd1 _02527_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09937__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ cpu.RF0.registers\[19\]\[11\] net616 net583 cpu.RF0.registers\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07412__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ net971 cpu.RF0.registers\[15\]\[14\] net829 vssd1 vssd1 vccd1 vccd1 _02389_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14261__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13829__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_2
Xfanout221 net223 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout232 net235 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 net267 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 _05846_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 _05688_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09808_ _03145_ net434 net289 _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__o211a_1
XANTENNA__10630__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _04392_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07505__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _05018_ _05025_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or3_4
XANTENNA__13979__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ net1466 net497 net280 cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07224__B cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ net2444 net251 net347 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ cpu.LCD0.row_2\[83\] net1755 net998 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13209__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ clknet_leaf_16_clk _01531_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11632_ net506 _05765_ _05907_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__and3_4
XANTENNA__12224__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__D1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07240__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ clknet_leaf_57_clk _01464_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11563_ net2699 net143 net369 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ clknet_leaf_31_clk cpu.RU0.next_FetchedData\[9\] net1206 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[9\] sky130_fd_sc_hd__dfrtp_1
X_10514_ net1135 a1.ADR_I\[1\] net915 _05644_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14282_ clknet_leaf_100_clk _01395_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13359__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11494_ net2062 net155 net374 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14604__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ clknet_leaf_44_clk _00413_ net1312 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09928__A1 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ net13 net754 net564 a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13164_ clknet_leaf_35_clk _00344_ net1259 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07403__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ cpu.f0.i\[0\] net270 vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ _05987_ _05995_ net557 vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__and3_4
XFILLER_0_23_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13095_ clknet_leaf_46_clk _00275_ net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_12046_ cpu.LCD0.cnt_500hz\[0\] cpu.LCD0.cnt_500hz\[1\] cpu.LCD0.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a21o_1
XANTENNA__08364__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11636__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13997_ clknet_leaf_102_clk _01110_ net1215 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_20_clk _00137_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10474__B2 a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12879_ clknet_leaf_1_clk cpu.c0.next_count\[10\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11371__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14134__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14618_ clknet_leaf_31_clk _01719_ net1208 vssd1 vssd1 vccd1 vccd1 cpu.f0.read_i
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12215__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A1 cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14549_ clknet_leaf_49_clk _01651_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10777__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ cpu.RF0.registers\[22\]\[25\] net670 _03345_ _03347_ _03350_ vssd1 vssd1
+ vccd1 vccd1 _03361_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload101 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_6
XANTENNA__14284__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07021_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09348__Y _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ cpu.RF0.registers\[5\]\[26\] net702 net665 _04251_ _04254_ vssd1 vssd1 vccd1
+ vccd1 _04263_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10016__A cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14486__RESET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ net1029 cpu.RF0.registers\[21\]\[30\] net795 vssd1 vssd1 vccd1 vccd1 _03214_
+ sky130_fd_sc_hd__and3_1
Xhold18 _01476_ vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 cpu.f0.data_adr\[19\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14415__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__B _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ net523 _03142_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_97_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12939__Q a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ cpu.CU0.funct3\[1\] cpu.CU0.funct3\[0\] cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1
+ vccd1 _02096_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06867__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07325__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07785_ _03061_ _03066_ _03067_ _03068_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__or4_1
XANTENNA__08107__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_A _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09524_ _02507_ _03698_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06736_ net936 cpu.RF0.registers\[10\]\[30\] net860 vssd1 vssd1 vccd1 vccd1 _02027_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09455_ _02982_ _04158_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06667_ a1.CPU_DAT_O\[3\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1273_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08406_ cpu.RF0.registers\[0\]\[10\] net664 net550 vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09607__B1 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09386_ net470 _04567_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07698__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06598_ _01970_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__inv_2
XANTENNA__14627__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07060__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ cpu.RF0.registers\[0\]\[12\] net661 net548 vssd1 vssd1 vccd1 vccd1 _03628_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07094__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ cpu.RF0.registers\[29\]\[15\] net673 _03556_ _03557_ _03558_ vssd1 vssd1
+ vccd1 vccd1 _03559_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07219_ net956 cpu.RF0.registers\[1\]\[9\] net804 vssd1 vssd1 vccd1 vccd1 _02510_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10625__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ cpu.RF0.registers\[10\]\[21\] net691 net684 cpu.RF0.registers\[24\]\[21\]
+ _03485_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a221o_1
XANTENNA__13651__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ cpu.f0.i\[7\] cpu.f0.i\[8\] net527 vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08322__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ cpu.IM0.address_IM\[27\] _05422_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1005 net1011 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_2
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14007__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1038 net1041 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11456__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
XANTENNA__09434__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ clknet_leaf_5_clk _01033_ net1148 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07235__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13851_ clknet_leaf_13_clk _00964_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14157__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ net2731 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__clkbuf_1
X_13782_ clknet_leaf_59_clk _00895_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ net988 cpu.f0.write_data\[20\] vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__or2_2
X_12733_ cpu.f0.i\[0\] _01872_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__or2_1
XANTENNA__11191__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12664_ net2828 net2585 net1001 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__mux2_1
XANTENNA__07872__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14403_ clknet_leaf_16_clk _01514_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.CU0.bit30
+ sky130_fd_sc_hd__dfrtp_4
X_11615_ net2829 net173 net361 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XANTENNA__09074__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ cpu.IM0.address_IM\[1\] _06353_ _06349_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__mux2_1
XANTENNA__07401__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ clknet_leaf_50_clk _01447_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfxtp_1
X_11546_ net2117 net208 net367 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14265_ clknet_leaf_42_clk _01378_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11477_ net2758 net217 net374 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
X_13216_ clknet_leaf_74_clk _00396_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ cpu.f0.i\[26\] net269 vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__nand2_1
XANTENNA__12899__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14196_ clknet_leaf_69_clk _01309_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07388__A1 cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07388__B2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13147_ clknet_leaf_53_clk _00327_ net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ cpu.f0.data_adr\[29\] net726 _05479_ _05592_ vssd1 vssd1 vccd1 vccd1 _00082_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09184__X _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13078_ clknet_leaf_53_clk _00258_ net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08337__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ cpu.LCD0.cnt_20ms\[2\] cpu.LCD0.cnt_20ms\[1\] cpu.LCD0.cnt_20ms\[0\] vssd1
+ vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07570_ _02857_ _02858_ _02859_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__or4_1
XANTENNA__09837__B1 _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06521_ cpu.f0.num\[21\] cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13524__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__B2 a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10998__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ _04422_ _04433_ net450 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__mux2_1
X_06452_ net2846 _01840_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07863__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ _04459_ _04461_ _02756_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
X_06383_ cpu.f0.num\[10\] vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13674__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ net1078 cpu.RF0.registers\[24\]\[23\] net870 vssd1 vssd1 vccd1 vccd1 _03413_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09359__X _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload51_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08053_ net939 cpu.RF0.registers\[6\]\[25\] net852 vssd1 vssd1 vccd1 vccd1 _03344_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07004_ net1034 cpu.RF0.registers\[27\]\[23\] net775 vssd1 vssd1 vccd1 vccd1 _02295_
+ sky130_fd_sc_hd__and3_1
Xmax_cap741 _01852_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09222__D1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08576__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__A1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__B2 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _04243_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__nor2_1
XANTENNA__07981__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13054__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06878__B net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _02213_ _03149_ _03172_ net488 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a31o_1
XANTENNA_hold1227_A cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ net934 cpu.RF0.registers\[15\]\[17\] net859 vssd1 vssd1 vccd1 vccd1 _04177_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10135__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ cpu.RF0.registers\[26\]\[24\] net600 net565 cpu.RF0.registers\[30\]\[24\]
+ _03127_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a221o_1
XANTENNA__10968__X _05863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07768_ net1042 cpu.RF0.registers\[22\]\[21\] net801 vssd1 vssd1 vccd1 vccd1 _03059_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08438__X _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _04737_ _04797_ net471 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06719_ net1114 net1116 net1110 net1112 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__nor4b_2
XANTENNA_fanout913_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ net1028 cpu.RF0.registers\[26\]\[17\] net786 vssd1 vssd1 vccd1 vccd1 _02990_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07303__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08500__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10989__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ _04535_ _04677_ _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__A2 _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08317__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ net478 _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__o21ai_1
X_11400_ net2201 net131 net386 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07606__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ net1119 net1694 net529 net1067 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08614__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11331_ net2442 net146 net396 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
X_14050_ clknet_leaf_10_clk _01163_ net1222 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11262_ net1873 net157 net402 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__mux2_1
XANTENNA__08901__X _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ clknet_leaf_36_clk _00190_ net1263 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08052__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _05472_ _05473_ _05474_ net126 net628 vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a221o_1
XANTENNA__08031__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ net2931 net153 net410 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ cpu.IM0.address_IM\[24\] _05387_ cpu.IM0.address_IM\[25\] vssd1 vssd1 vccd1
+ vccd1 _05412_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11186__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__inv_2
X_13903_ clknet_leaf_87_clk _01016_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13547__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__X _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11914__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13834_ clknet_leaf_99_clk _00947_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09180__A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__X _02543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13765_ clknet_leaf_10_clk _00878_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ net1883 net928 net276 _05869_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a22o_1
XANTENNA__08098__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09295__A1 _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13697__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12716_ net2238 cpu.LCD0.row_2\[110\] net1006 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__mux2_1
XANTENNA__06803__C_N cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13696_ clknet_leaf_9_clk _00809_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ net2691 net2499 net1009 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07058__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _06341_ cpu.SR1.char_in\[4\] _06320_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08524__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__B1 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14317_ clknet_leaf_103_clk _01430_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ net2057 net145 net372 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__mux2_1
XANTENNA__08270__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 cpu.RF0.registers\[23\]\[30\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold318 cpu.RF0.registers\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12854__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14248_ clknet_leaf_98_clk _01361_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold329 cpu.RF0.registers\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12354__A1 cpu.K0.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13077__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__C1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14179_ clknet_leaf_77_clk _01292_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14322__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07574__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _04029_ _04030_ _03934_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__a21o_1
Xhold1007 cpu.RF0.registers\[10\]\[18\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1018 cpu.RF0.registers\[28\]\[10\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1029 cpu.RF0.registers\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1380 net1384 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14472__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08671_ _03951_ _03956_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or3_4
XANTENNA__13027__D net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11824__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ net960 cpu.RF0.registers\[12\]\[13\] net765 vssd1 vssd1 vccd1 vccd1 _02913_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12914__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12409__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload99_A clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12866__D net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07553_ net969 cpu.RF0.registers\[6\]\[8\] net803 vssd1 vssd1 vccd1 vccd1 _02844_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09286__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ _01780_ cpu.f0.state\[3\] net528 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a21o_1
XANTENNA__07297__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12290__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07836__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ net1060 cpu.RF0.registers\[28\]\[5\] net767 vssd1 vssd1 vccd1 vccd1 _02775_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _04414_ _04478_ _04495_ net302 _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a221o_1
X_06435_ _01829_ _01833_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07041__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout327_A _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__X _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09154_ _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__nor2_2
X_06366_ net1071 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08105_ cpu.RF0.registers\[1\]\[22\] net714 net674 cpu.RF0.registers\[6\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09994__C1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09085_ net495 net460 net454 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__and3_1
XANTENNA__08261__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08036_ cpu.RF0.registers\[28\]\[24\] net706 _03306_ _03313_ _03318_ vssd1 vssd1
+ vccd1 vccd1 _03327_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_13_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold830 _00330_ vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold841 cpu.LCD0.row_2\[98\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold852 cpu.RF0.registers\[16\]\[18\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__C1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 cpu.RF0.registers\[8\]\[23\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 cpu.LCD0.row_2\[64\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold885 cpu.LCD0.row_2\[18\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold896 cpu.RF0.registers\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ cpu.IM0.address_IM\[13\] _02904_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08938_ cpu.RF0.registers\[3\]\[27\] net645 net640 cpu.RF0.registers\[19\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__a22o_1
Xhold1530 a1.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1 net2936 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ net490 _02945_ _02983_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_4_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net2554 net183 net431 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
XANTENNA__09712__B _04405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ net2924 net205 net326 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08609__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ net2003 net236 net432 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13312__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ clknet_leaf_4_clk _00663_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12281__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ cpu.f0.data_adr\[14\] _05086_ net990 vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ _05534_ _06267_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ clknet_leaf_105_clk _00594_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12565__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ cpu.LCD0.row_1\[99\] net2623 net898 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
X_12432_ net2903 net534 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12862__Q cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__B2 _06345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ net1122 net1434 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10595__A0 cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14345__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14102_ clknet_leaf_58_clk _01215_ net1367 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11314_ net1751 net201 net395 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__mux2_1
X_12294_ cpu.LCD0.row_1\[87\] _05986_ _06105_ _06157_ _06187_ vssd1 vssd1 vccd1 vccd1
+ _06188_ sky130_fd_sc_hd__a2111o_1
X_14033_ clknet_leaf_77_clk _01146_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11909__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ net2067 net217 net402 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08004__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14100__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07212__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10898__A1 _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ net2721 net230 net412 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__mux2_1
XANTENNA__14495__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05361_ _05372_ _05393_ _02310_ cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1
+ vccd1 _05396_ sky130_fd_sc_hd__a32o_1
XANTENNA__12937__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10058_ net127 _05332_ _05331_ net630 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__a211o_1
XANTENNA__07126__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09622__B _03233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08078__X _03369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13817_ clknet_leaf_91_clk _00930_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09268__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12272__B1 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_72_clk _00861_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ clknet_leaf_87_clk _00792_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08491__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07796__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 _00178_ vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _00167_ vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 net81 vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13712__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 cpu.RF0.registers\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11819__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 cpu.RF0.registers\[0\]\[9\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _05183_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nand2_1
Xhold159 cpu.RF0.registers\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout606 _02144_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09841_ _03540_ _05076_ _03538_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a21oi_1
Xfanout617 net620 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09085__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09743__A2 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06502__A cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_2
Xfanout639 _02065_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
XANTENNA_clkload14_A clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08951__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ net486 _04758_ _05062_ _04410_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13862__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06984_ net544 _02271_ _02273_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09372__X _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ cpu.RF0.registers\[15\]\[0\] net946 net857 vssd1 vssd1 vccd1 vccd1 _04014_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07036__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09091__Y _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ net1102 cpu.RF0.registers\[19\]\[2\] _02062_ vssd1 vssd1 vccd1 vccd1 _03945_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10510__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14218__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06875__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07605_ cpu.RF0.registers\[23\]\[12\] net614 _02879_ _02884_ _02886_ vssd1 vssd1
+ vccd1 vccd1 _02896_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07333__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ net1100 cpu.RF0.registers\[28\]\[4\] net868 vssd1 vssd1 vccd1 vccd1 _03876_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09259__B2 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07536_ cpu.RF0.registers\[15\]\[6\] _02167_ _02826_ net622 vssd1 vssd1 vccd1 vccd1
+ _02827_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07467_ net487 net476 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_27_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13242__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14368__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ net306 _04409_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06418_ cpu.c0.count\[5\] cpu.c0.count\[6\] cpu.c0.count\[7\] cpu.c0.count\[4\] vssd1
+ vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__or4bb_1
X_07398_ net971 cpu.RF0.registers\[5\]\[0\] net797 vssd1 vssd1 vccd1 vccd1 _02689_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08164__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09137_ net462 _03866_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nor2_1
XANTENNA__10577__A0 cpu.f0.write_data\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_X net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09068_ net438 _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__or2_1
XANTENNA__13392__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ net947 cpu.RF0.registers\[11\]\[24\] net879 vssd1 vssd1 vccd1 vccd1 _03310_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10633__S net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 cpu.RF0.registers\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 a1.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 cpu.RF0.registers\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ cpu.IG0.Instr\[7\] cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__nor2_2
Xhold693 cpu.RF0.registers\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14402__Q cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07942__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_44_clk net1426 net1305 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10869__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11464__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1360 cpu.RF0.registers\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 cpu.RF0.registers\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1382 cpu.RF0.registers\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ net2342 net249 net321 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
XANTENNA__10501__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1393 cpu.f0.num\[5\] vssd1 vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08339__A _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14651_ clknet_leaf_22_clk _01752_ net1172 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11863_ net505 _05912_ _05920_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__and3_4
XFILLER_0_32_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10814_ cpu.f0.data_adr\[29\] _04551_ net991 vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__mux2_1
X_13602_ clknet_leaf_102_clk _00715_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14582_ clknet_leaf_47_clk _01684_ net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_11794_ net2309 net142 net341 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10804__A1 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10745_ cpu.IM0.address_IM\[9\] net1017 _05688_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_
+ sky130_fd_sc_hd__a22o_1
X_13533_ clknet_leaf_66_clk _00646_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13464_ clknet_leaf_6_clk _00577_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ net2564 cpu.LCD0.row_1\[90\] net897 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13735__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12415_ net1512 net732 net501 _06231_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__o22a_1
XANTENNA__08225__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ clknet_leaf_68_clk _00508_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12346_ cpu.LCD0.cnt_20ms\[15\] _06213_ net1368 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08802__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06787__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11639__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net1370 _06170_ _06171_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13885__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ clknet_leaf_5_clk _01129_ net1145 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07418__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ net1962 net159 net407 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ net1815 net165 net417 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13115__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09633__A _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10779__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11374__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13265__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__B1 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ cpu.RF0.registers\[5\]\[11\] net702 net666 _03659_ _03660_ vssd1 vssd1 vccd1
+ vccd1 _03661_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07321_ net1062 cpu.RF0.registers\[16\]\[3\] net832 vssd1 vssd1 vccd1 vccd1 _02612_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ cpu.RF0.registers\[0\]\[9\] net617 _02539_ _02542_ vssd1 vssd1 vccd1 vccd1
+ _02543_ sky130_fd_sc_hd__o22a_2
XFILLER_0_27_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08415__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ cpu.CU0.bit30 net520 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09413__B2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11549__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12234__A _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07328__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A2 _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout403 _05919_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_4
Xfanout414 net417 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout425 _05913_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_8
Xfanout436 _04403_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_A _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _05109_ _05110_ _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__or3_2
Xfanout447 _03300_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1101_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout469 _02717_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
X_09755_ net450 _04435_ _04437_ _05045_ _02758_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__o311a_1
X_06967_ cpu.RF0.registers\[13\]\[25\] net597 net588 cpu.RF0.registers\[1\]\[25\]
+ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06886__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ cpu.RF0.registers\[20\]\[0\] net709 net641 cpu.RF0.registers\[19\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a22o_1
XANTENNA__11287__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09686_ _04975_ _04976_ _04974_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a21oi_1
X_06898_ net966 net766 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ cpu.RF0.registers\[3\]\[3\] net643 _03926_ _03927_ net668 vssd1 vssd1 vccd1
+ vccd1 _03928_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_29_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1091_X net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__B cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08568_ cpu.RF0.registers\[11\]\[5\] net688 net683 cpu.RF0.registers\[15\]\[5\] _03840_
+ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07350__X _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ net978 cpu.RF0.registers\[13\]\[6\] net794 vssd1 vssd1 vccd1 vccd1 _02810_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ cpu.RF0.registers\[5\]\[7\] net703 net688 cpu.RF0.registers\[11\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1356_X net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10530_ net1132 net2409 net912 _05652_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_94_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire815 _02137_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ net10 net754 net564 a1.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__a22o_1
XANTENNA__08207__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ cpu.LCD0.row_2\[115\] _06007_ _06021_ cpu.LCD0.row_1\[91\] vssd1 vssd1 vccd1
+ vccd1 _06098_ sky130_fd_sc_hd__a22o_1
X_13180_ clknet_leaf_30_clk _00360_ net1207 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ cpu.f0.i\[8\] net271 vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ cpu.LCD0.row_1\[40\] _06030_ _06031_ cpu.LCD0.row_1\[24\] _06029_ vssd1 vssd1
+ vccd1 vccd1 _06032_ sky130_fd_sc_hd__a221o_1
XANTENNA__11459__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ _05969_ net502 _05968_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__and3b_1
Xhold490 cpu.RF0.registers\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08060__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ cpu.f0.write_data\[26\] _05894_ net985 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__mux2_1
XANTENNA__10722__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net984 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_2
Xfanout992 net994 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11194__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13288__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12964_ clknet_leaf_44_clk net1517 net1305 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XANTENNA__14533__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1190 cpu.RF0.registers\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11915_ net2481 net185 net323 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
XANTENNA__07404__C net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__X _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ clknet_leaf_28_clk _00009_ net1188 vssd1 vssd1 vccd1 vccd1 a1.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08694__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634_ clknet_leaf_31_clk _01735_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ net1922 net173 net332 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07701__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14565_ clknet_leaf_47_clk _01667_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_11777_ net2068 net209 net339 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__mux2_1
XANTENNA__08446__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10789__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10728_ cpu.IM0.address_IM\[4\] net1015 net285 _05695_ vssd1 vssd1 vccd1 vccd1 _05696_
+ sky130_fd_sc_hd__a22o_1
X_13516_ clknet_leaf_79_clk _00629_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14496_ clknet_leaf_35_clk _01598_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_77_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10659_ net2907 net2737 net906 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
X_13447_ clknet_leaf_81_clk _00560_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload13 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload24 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinv_2
Xclkload35 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinv_8
Xclkload46 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload46/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09628__A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09946__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_94_clk _00491_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload57 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_24_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload68 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10556__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload79 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_8
X_12329_ _06203_ _06204_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__nor2_1
XANTENNA__12054__A _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B1 _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ cpu.RF0.registers\[26\]\[28\] net600 net597 cpu.RF0.registers\[13\]\[28\]
+ _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__a221o_1
X_06821_ cpu.CU0.funct3\[2\] _02103_ _02107_ _02097_ vssd1 vssd1 vccd1 vccd1 _02112_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_78_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _03769_ _04040_ _03735_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21oi_1
X_06752_ net1081 cpu.RF0.registers\[29\]\[30\] net848 vssd1 vssd1 vccd1 vccd1 _02043_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09331__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ _04720_ _04761_ net472 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13900__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06683_ a1.CPU_DAT_O\[19\] net889 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[19\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08685__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11832__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08422_ net936 cpu.RF0.registers\[2\]\[9\] net855 vssd1 vssd1 vccd1 vccd1 _03713_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12218__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07893__B1 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ net1093 cpu.RF0.registers\[27\]\[11\] net879 vssd1 vssd1 vccd1 vccd1 _03644_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12769__B2 cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout142_A _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07304_ cpu.RF0.registers\[9\]\[4\] net573 net568 cpu.RF0.registers\[25\]\[4\] _02594_
+ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a221o_1
XANTENNA__11441__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ net1082 cpu.RF0.registers\[16\]\[13\] net841 vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload7 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
X_07235_ net959 cpu.RF0.registers\[9\]\[9\] net758 vssd1 vssd1 vccd1 vccd1 _02526_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_73_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ net969 cpu.RF0.registers\[8\]\[11\] net812 vssd1 vssd1 vccd1 vccd1 _02457_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08442__A _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07984__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14406__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11279__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07097_ net1049 cpu.RF0.registers\[28\]\[14\] net767 vssd1 vssd1 vccd1 vccd1 _02388_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1316_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout200 _05802_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
Xfanout1209 net1210 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 _05799_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold1424_A cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10911__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout244 _05778_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13430__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14556__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06897__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A1 cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09273__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _04695_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
X_09807_ net294 net297 _04917_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__mux2_1
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 _04392_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
X_07999_ cpu.RF0.registers\[27\]\[28\] net711 _03272_ _03278_ _03280_ vssd1 vssd1
+ vccd1 vccd1 _03290_ sky130_fd_sc_hd__a2111o_1
X_09738_ net471 _04440_ _04564_ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10212__A cpu.IM0.address_IM\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13580__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ _04949_ _04959_ _04958_ _04957_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o211a_1
XANTENNA__07224__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11700_ net2519 net253 net348 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10483__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ net2483 cpu.LCD0.row_2\[74\] net1001 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XANTENNA__07884__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11631_ net2742 net130 net358 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08428__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14350_ clknet_leaf_28_clk _01463_ net1185 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11562_ net2181 net146 net368 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ net51 net917 vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__and2_1
X_13301_ clknet_leaf_31_clk cpu.RU0.next_FetchedData\[8\] net1205 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08055__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14281_ clknet_leaf_105_clk _01394_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11493_ net1907 net159 net375 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13232_ clknet_leaf_44_clk _00412_ net1312 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ net2 net753 net562 a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__o22a_1
XANTENNA__09928__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14086__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10538__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13163_ clknet_leaf_53_clk net1581 net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10375_ _01939_ _05477_ _05601_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__or3_1
XANTENNA__09167__B _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08600__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__B1 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net746 _05993_ _05996_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and3_4
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13094_ clknet_leaf_53_clk net2217 net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_clk_X clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ _01953_ _05957_ _05959_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07167__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13923__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ clknet_leaf_74_clk _01109_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12808__RESET_B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_20_clk _00136_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08667__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11652__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12878_ clknet_leaf_0_clk cpu.c0.next_count\[9\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[9\] sky130_fd_sc_hd__dfrtp_1
X_14617_ clknet_leaf_33_clk cpu.f0.next_lcd_en net1247 vssd1 vssd1 vccd1 vccd1 cpu.SR1.enable
+ sky130_fd_sc_hd__dfrtp_1
X_11829_ net1943 net131 net334 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14548_ clknet_leaf_46_clk net2339 net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13303__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14429__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14479_ clknet_leaf_30_clk _00005_ net1208 vssd1 vssd1 vccd1 vccd1 cpu.RU0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload102 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_12
X_07020_ _02309_ _02310_ net522 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_4
XFILLER_0_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09358__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11099__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13453__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14579__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ _04248_ _04255_ _04260_ _04261_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__or4_1
XANTENNA__11827__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ net1030 cpu.RF0.registers\[16\]\[30\] net831 vssd1 vssd1 vccd1 vccd1 _03213_
+ sky130_fd_sc_hd__and3_1
Xhold19 a1.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A2 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ net544 _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06804_ cpu.CU0.funct3\[2\] cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__nor2_1
X_07784_ cpu.RF0.registers\[7\]\[21\] net596 _03074_ net624 vssd1 vssd1 vccd1 vccd1
+ _03075_ sky130_fd_sc_hd__a211o_1
XANTENNA__10032__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ _03735_ _04040_ _04043_ _04045_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__o211ai_2
X_06735_ net944 net861 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__and2_1
XANTENNA__11562__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _05932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__Y _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _02982_ _04158_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1099_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06666_ a1.CPU_DAT_O\[2\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07866__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10465__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08405_ _03685_ _03688_ _03692_ _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__or4_1
XANTENNA__12955__Q a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _02348_ _04402_ net291 _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a211o_1
XANTENNA__09607__A1 _04025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06597_ net1366 _01969_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout524_A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _03617_ _03618_ _03623_ _03626_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07094__A1 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__Y _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ cpu.RF0.registers\[8\]\[15\] net707 net681 cpu.RF0.registers\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ cpu.IG0.Instr\[29\] net522 net520 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__and3_1
X_08198_ cpu.RF0.registers\[28\]\[21\] net705 _03478_ _03481_ _03487_ vssd1 vssd1
+ vccd1 vccd1 _03489_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout893_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07149_ net966 cpu.RF0.registers\[1\]\[11\] net805 vssd1 vssd1 vccd1 vccd1 _02440_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08043__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10160_ cpu.IM0.address_IM\[26\] net932 _05425_ _05426_ vssd1 vssd1 vccd1 vccd1 _00049_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13946__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1006 net1011 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11737__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1017 cpu.RU0.state\[5\] vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
XANTENNA__10641__S net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ cpu.IM0.address_IM\[20\] _03042_ _05352_ vssd1 vssd1 vccd1 vccd1 _05363_
+ sky130_fd_sc_hd__a21o_1
Xfanout1028 net1033 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_2
Xfanout1039 net1041 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09207__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12141__B _01965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12970__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ clknet_leaf_94_clk _00963_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ net2633 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__clkbuf_1
X_10993_ net282 _05880_ net995 vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__o21ai_1
X_13781_ clknet_leaf_73_clk _00894_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09846__B2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11472__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ cpu.f0.state\[7\] net499 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08347__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_52_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12663_ net2524 cpu.LCD0.row_2\[57\] net1009 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14402_ clknet_leaf_23_clk _01513_ net1194 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12602__A0 cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10208__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ net2682 net195 net360 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12594_ _05058_ _06352_ net625 vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14333_ clknet_leaf_56_clk _01446_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11545_ net2825 net204 net367 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XANTENNA__13476__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08821__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_67_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14264_ clknet_leaf_8_clk _01377_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11476_ net1703 net222 net376 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08513__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11995__X _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net1125 _05631_ net264 net2211 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__a2bb2o_1
X_13215_ clknet_leaf_95_clk _00395_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14195_ clknet_leaf_68_clk _01308_ net1324 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10117__A cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07388__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ clknet_leaf_52_clk net2430 net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_10358_ net528 _05588_ _05591_ net308 vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a22o_1
XANTENNA__11647__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ clknet_leaf_51_clk _00257_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09625__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _01810_ _05529_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ net2876 cpu.LCD0.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10144__A1 cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14101__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07560__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10787__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ clknet_leaf_94_clk _01092_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09837__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ cpu.f0.num\[22\] net1019 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nand2_1
XANTENNA__11235__X _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07799__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14251__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06451_ net1440 _01827_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[8\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13819__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09170_ net469 _03699_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a21oi_1
X_06382_ cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ net1076 cpu.RF0.registers\[17\]\[23\] net882 vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08273__B1 _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09088__A _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ net939 cpu.RF0.registers\[7\]\[25\] net847 vssd1 vssd1 vccd1 vccd1 _03343_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkload44_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12843__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ net1035 cpu.RF0.registers\[23\]\[23\] net816 vssd1 vssd1 vccd1 vccd1 _02294_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_24_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08423__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap742 _01850_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_2
XFILLER_0_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08576__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07379__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07039__C _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__Y _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _02213_ _03149_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1014_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__inv_2
XANTENNA__10135__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08885_ net935 cpu.RF0.registers\[5\]\[17\] net866 vssd1 vssd1 vccd1 vccd1 _04176_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout474_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ cpu.RF0.registers\[17\]\[24\] net606 net572 cpu.RF0.registers\[12\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13349__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net1042 cpu.RF0.registers\[17\]\[21\] net805 vssd1 vssd1 vccd1 vccd1 _03058_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout641_A _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _04795_ _04796_ net457 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07839__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06718_ net1090 net880 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__and2_1
XANTENNA__08167__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07698_ net1031 cpu.RF0.registers\[25\]\[17\] net756 vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07071__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ _03019_ net439 _04726_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__o22ai_1
X_06649_ a1.CPU_DAT_O\[17\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[17\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13499__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _04385_ _04524_ _04529_ net301 _04382_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09056__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08319_ net1086 cpu.RF0.registers\[21\]\[12\] net866 vssd1 vssd1 vccd1 vccd1 _03610_
+ sky130_fd_sc_hd__and3_1
X_09299_ _04367_ _04419_ net475 vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ net1821 net148 net394 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XANTENNA__10071__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ net1623 net160 net403 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13000_ clknet_leaf_36_clk _00189_ net1260 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09285__X _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ cpu.IM0.address_IM\[31\] _05464_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__xor2_1
XANTENNA__09764__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ net1958 net163 net410 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10143_ cpu.IM0.address_IM\[25\] cpu.IM0.address_IM\[24\] _05387_ vssd1 vssd1 vccd1
+ vccd1 _05411_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10224__X _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12449__B1_N net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input35_A gpio_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10074_ cpu.IM0.address_IM\[18\] _02349_ _05336_ _05335_ vssd1 vssd1 vccd1 vccd1
+ _05347_ sky130_fd_sc_hd__a31o_1
XANTENNA__10126__A1 _05328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13902_ clknet_leaf_1_clk _01015_ net1139 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14274__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ clknet_leaf_103_clk _00946_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09180__B _04025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13764_ clknet_leaf_96_clk _00877_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10976_ net991 cpu.f0.write_data\[15\] _05852_ _05867_ vssd1 vssd1 vccd1 vccd1 _05869_
+ sky130_fd_sc_hd__o22a_1
X_12715_ cpu.LCD0.row_2\[117\] cpu.LCD0.row_2\[109\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ clknet_leaf_106_clk _00808_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07845__A3 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ net2351 net2285 net1008 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08255__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ _06308_ _06337_ _06340_ net1128 vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06805__A1 cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14316_ clknet_leaf_68_clk _01429_ net1296 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11528_ net1775 net150 net370 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 cpu.RF0.registers\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 cpu.RF0.registers\[24\]\[17\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ clknet_leaf_81_clk _01360_ net1291 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11459_ net2562 net178 net380 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XANTENNA__10365__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_94_clk _01291_ net1227 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11377__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ clknet_leaf_48_clk _00309_ net1355 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[93\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07781__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07156__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 a1.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12823__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14617__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 cpu.RF0.registers\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14047__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1370 net1371 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__clkbuf_4
X_08670_ _03957_ _03958_ _03959_ _03960_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__or4_1
Xfanout1381 net1383 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07533__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net960 cpu.RF0.registers\[4\]\[13\] net780 vssd1 vssd1 vccd1 vccd1 _02912_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__B _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13641__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07552_ net1051 cpu.RF0.registers\[29\]\[8\] net793 vssd1 vssd1 vccd1 vccd1 _02843_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12001__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06503_ cpu.K0.keyvalid cpu.f0.state\[5\] _01890_ vssd1 vssd1 vccd1 vccd1 _01893_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08418__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07483_ net982 cpu.RF0.registers\[7\]\[5\] net818 vssd1 vssd1 vccd1 vccd1 _02774_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08494__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07322__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11840__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06434_ cpu.c0.count\[15\] _01842_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__and2_1
X_09222_ net478 _04504_ _04507_ _04512_ net278 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ net302 _04411_ _04414_ _04442_ _04408_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13791__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06365_ net1051 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08104_ cpu.RF0.registers\[5\]\[22\] net702 net680 cpu.RF0.registers\[18\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09084_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ cpu.RF0.registers\[26\]\[24\] net639 _03307_ _03308_ _03317_ vssd1 vssd1
+ vccd1 vccd1 _03326_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13021__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold820 cpu.LCD0.row_1\[32\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10980__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14147__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 cpu.RF0.registers\[1\]\[30\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 _01689_ vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 cpu.RF0.registers\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07992__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold864 a1.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold875 cpu.RF0.registers\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold886 cpu.RF0.registers\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold897 cpu.LCD0.row_1\[27\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ cpu.IM0.address_IM\[12\] net931 _05265_ _05266_ vssd1 vssd1 vccd1 vccd1 _00035_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13171__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14297__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ cpu.RF0.registers\[31\]\[27\] net687 net684 cpu.RF0.registers\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__a22o_1
XANTENNA__10108__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1520 cpu.LCD0.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1 net2926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 cpu.LCD0.row_1\[54\] vssd1 vssd1 vccd1 vccd1 net2937 sky130_fd_sc_hd__dlygate4sd3_1
X_08868_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _03106_ _03107_ _03108_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__or4_1
X_08799_ net441 _04088_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1386_X net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ _05768_ _05769_ cpu.IM0.address_IM\[0\] _02001_ vssd1 vssd1 vccd1 vccd1 _05770_
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_36_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ net1913 net561 net539 _05719_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__a22o_1
XANTENNA__12281__A1 cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07232__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ net1021 _05526_ net257 cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__a31o_1
X_10692_ net2311 net2235 net897 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
X_13480_ clknet_leaf_97_clk _00593_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08237__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ net1740 net731 net501 _06239_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12584__A2 cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ net1122 net1566 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and2_1
XANTENNA__08063__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ clknet_leaf_73_clk _01214_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11313_ net2079 net212 net395 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__mux2_1
X_12293_ cpu.LCD0.row_2\[111\] _06012_ _06028_ cpu.LCD0.row_1\[119\] vssd1 vssd1 vccd1
+ vccd1 _06187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09737__B1 _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09456__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ clknet_leaf_75_clk _01145_ net1334 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11244_ net1714 net220 net404 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13514__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11197__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07212__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ net1777 net232 net412 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__mux2_1
X_10126_ _05328_ _05348_ _05350_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11925__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__Y _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13664__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ cpu.IM0.address_IM\[18\] _05319_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__xor2_1
XANTENNA__07704__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload0_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13816_ clknet_leaf_6_clk _00929_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09268__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13747_ clknet_leaf_69_clk _00860_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10959_ _02506_ net516 _05852_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11660__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10283__B1 cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10822__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13678_ clknet_leaf_4_clk _00791_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ cpu.LCD0.row_2\[31\] net2465 net1004 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08228__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09976__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 cpu.RF0.registers\[0\]\[11\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 cpu.FetchedInstr\[13\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold127 cpu.FetchedInstr\[28\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net87 vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14299__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09840_ net512 _05122_ _05123_ net258 _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__o311a_2
Xfanout607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_8
Xfanout629 net632 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
XANTENNA__06557__A3 _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08951__A1 cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ net474 _04522_ net485 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07317__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06983_ net544 _02271_ _02273_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a21o_1
XANTENNA__06962__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11835__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ cpu.RF0.registers\[6\]\[0\] net675 net667 _04011_ _04012_ vssd1 vssd1 vccd1
+ vccd1 _04013_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_33_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__A1 _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net1102 cpu.RF0.registers\[27\]\[2\] net879 vssd1 vssd1 vccd1 vccd1 _03944_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_53_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout172_A _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07604_ cpu.RF0.registers\[10\]\[12\] net569 _02878_ _02882_ _02889_ vssd1 vssd1
+ vccd1 vccd1 _02895_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08584_ net1100 cpu.RF0.registers\[29\]\[4\] net849 vssd1 vssd1 vccd1 vccd1 _03875_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07901__X _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07535_ cpu.RF0.registers\[20\]\[6\] net594 net567 cpu.RF0.registers\[11\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1081_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout437_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07466_ net523 _02754_ _02755_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07987__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ net306 _04409_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nor2_2
X_06417_ cpu.c0.count\[13\] cpu.c0.count\[12\] cpu.c0.count\[14\] cpu.c0.count\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__or4b_1
XANTENNA__07690__A1 cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ net1048 cpu.RF0.registers\[23\]\[0\] net818 vssd1 vssd1 vccd1 vccd1 _02688_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout604_A _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1346_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09136_ _04419_ _04426_ net475 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10577__A1 _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__X _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13537__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09067_ cpu.IG0.Instr\[31\] _04357_ net543 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_92_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10914__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__A0 _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09276__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ net1099 cpu.RF0.registers\[31\]\[24\] net857 vssd1 vssd1 vccd1 vccd1 _03309_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07993__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 cpu.RF0.registers\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 cpu.RF0.registers\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12414__B _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 cpu.RF0.registers\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold683 cpu.RF0.registers\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 cpu.RF0.registers\[1\]\[23\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13687__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _05235_ _05238_ _05234_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ clknet_leaf_28_clk _00169_ net1188 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_71_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12430__A cpu.DM0.data_i\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10869__B _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1350 cpu.RF0.registers\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 cpu.LCD0.row_1\[64\] vssd1 vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07524__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11931_ net2558 net256 net321 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
Xhold1372 cpu.RF0.registers\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1383 cpu.LCD0.row_2\[57\] vssd1 vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__B2 a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1394 cpu.RF0.registers\[8\]\[8\] vssd1 vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
X_14650_ clknet_leaf_22_clk _01751_ net1173 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11862_ net2228 net131 net330 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ clknet_leaf_64_clk _00714_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ net1745 net561 net537 _05756_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__a22o_1
X_14581_ clknet_leaf_49_clk _01683_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[92\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__13067__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11793_ net2242 net147 net340 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11480__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ clknet_leaf_15_clk _00645_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ cpu.f0.data_adr\[9\] _04846_ net990 vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__mux2_1
XANTENNA__08355__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13463_ clknet_leaf_64_clk _00576_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ net2607 net2508 net906 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_80_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ cpu.DM0.data_i\[15\] _05847_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and2_1
X_13394_ clknet_leaf_69_clk _00507_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14462__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12345_ _06213_ _06214_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12904__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14392__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12276_ net111 net555 vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08090__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ clknet_leaf_0_clk _01128_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08521__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ net2058 net178 net408 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
XANTENNA__12190__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__X _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11158_ net2275 net169 net417 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11655__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10109_ net627 _04617_ net930 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a21oi_1
X_11089_ net2343 net170 net425 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XANTENNA__09633__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10779__B _04683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07434__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__A1_N _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11390__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ net974 cpu.RF0.registers\[11\]\[3\] net777 vssd1 vssd1 vccd1 vccd1 _02611_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09661__A2 _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07251_ _02533_ _02534_ _02540_ _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07182_ net546 _02470_ _02438_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a21o_2
XFILLER_0_26_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire774_A _02172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10734__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08271__Y _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__Y _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout404 _05919_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07727__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 _05911_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_6
X_09823_ _04566_ _04629_ _04634_ net272 _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__a221o_1
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout448 _03268_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 _02756_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10192__C1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net450 _05020_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__nand2_1
X_06966_ cpu.RF0.registers\[7\]\[25\] net595 net586 cpu.RF0.registers\[4\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a22o_1
XANTENNA__12958__Q a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ _03993_ _03994_ _03992_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ net476 _03964_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nand2_1
XANTENNA__08688__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ net963 cpu.RF0.registers\[9\]\[27\] net757 vssd1 vssd1 vccd1 vccd1 _02188_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout554_A _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1296_A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14335__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ cpu.RF0.registers\[1\]\[3\] _02007_ _03906_ _03908_ _03912_ vssd1 vssd1 vccd1
+ vccd1 _03927_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_16_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10201__C _05443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12396__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _03854_ _03855_ _03856_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ net1057 cpu.RF0.registers\[25\]\[6\] net759 vssd1 vssd1 vccd1 vccd1 _02809_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10798__A1 cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07112__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ cpu.RF0.registers\[20\]\[7\] net709 net707 cpu.RF0.registers\[8\]\[7\] _03779_
+ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ net976 cpu.RF0.registers\[13\]\[1\] net794 vssd1 vssd1 vccd1 vccd1 _02740_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07510__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08860__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12927__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10460_ net9 net752 net562 net2270 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__inv_2
X_10391_ net1125 _05613_ net264 net2155 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12130_ net745 _05981_ _05984_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and3_4
XANTENNA__07966__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07820__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ cpu.LCD0.cnt_500hz\[7\] cpu.LCD0.cnt_500hz\[8\] _05966_ vssd1 vssd1 vccd1
+ vccd1 _05969_ sky130_fd_sc_hd__and3_1
Xhold480 cpu.RF0.registers\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold491 cpu.LCD0.row_2\[103\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__B1 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11012_ _02247_ net532 net282 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06710__X _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A1 cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_2
Xfanout971 net973 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07254__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12868__Q cpu.K0.enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ clknet_leaf_44_clk net1459 net1305 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_84_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 cpu.RF0.registers\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 cpu.RF0.registers\[14\]\[24\] vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ net1699 net192 net322 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ clknet_leaf_28_clk _00008_ net1183 vssd1 vssd1 vccd1 vccd1 a1.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07541__X _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633_ clknet_leaf_26_clk _01734_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13702__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ net2733 net195 net332 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ clknet_leaf_47_clk _01666_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08085__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11776_ net1565 net204 net339 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__mux2_1
XANTENNA__07103__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08516__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13515_ clknet_leaf_91_clk _00628_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ cpu.f0.data_adr\[4\] _05016_ net994 vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14495_ clknet_leaf_33_clk _01597_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07420__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13852__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ clknet_leaf_6_clk _00559_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10658_ net2767 cpu.LCD0.row_1\[72\] net910 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08813__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload14 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_58_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload25 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08603__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload36 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_16
Xclkload47 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload47/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09946__A3 _05229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13377_ clknet_leaf_66_clk _00490_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09628__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10589_ cpu.f0.write_data\[6\] _02829_ net995 vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_16
XFILLER_0_2_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload69 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__clkinv_2
X_12328_ net2787 _06202_ net1340 vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10961__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ cpu.LCD0.row_2\[38\] _06004_ _06030_ cpu.LCD0.row_1\[46\] _06153_ vssd1 vssd1
+ vccd1 vccd1 _06154_ sky130_fd_sc_hd__a221o_1
XANTENNA__07148__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11385__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13232__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _02099_ _02106_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__nor3_1
X_06751_ net1088 net848 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__and2_2
XFILLER_0_56_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_75_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08134__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A1 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _04759_ _04760_ net457 vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06682_ net2816 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[18\] sky130_fd_sc_hd__and2_1
XFILLER_0_17_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13382__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08421_ net1078 cpu.RF0.registers\[21\]\[9\] net866 vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12769__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08352_ net1087 cpu.RF0.registers\[17\]\[11\] net883 vssd1 vssd1 vccd1 vccd1 _03643_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09095__A0 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ net1063 cpu.RF0.registers\[31\]\[4\] net829 net597 cpu.RF0.registers\[13\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08283_ net1086 cpu.RF0.registers\[29\]\[13\] net848 vssd1 vssd1 vccd1 vccd1 _03574_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07330__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07234_ net1035 cpu.RF0.registers\[20\]\[9\] net780 vssd1 vssd1 vccd1 vccd1 _02525_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_55_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07165_ net1043 cpu.RF0.registers\[23\]\[11\] net817 vssd1 vssd1 vccd1 vccd1 _02456_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1044_A cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07339__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07096_ cpu.RF0.registers\[24\]\[14\] net607 net584 cpu.RF0.registers\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1211_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12154__B1 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net204 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
Xfanout212 net215 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1309_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout223 _05788_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout671_A _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xfanout245 _05776_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XANTENNA__11295__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 _05772_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 _05605_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08373__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _03340_ _04204_ _04211_ net511 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a31o_1
XANTENNA__09570__B2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout278 _04382_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
X_07998_ cpu.RF0.registers\[8\]\[28\] net707 net675 cpu.RF0.registers\[6\]\[28\] _03288_
+ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a221o_1
XANTENNA__07074__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _05027_ _05026_ _03931_ net487 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__o2bb2a_1
X_06949_ cpu.RF0.registers\[8\]\[26\] net611 _02225_ _02227_ _02232_ vssd1 vssd1 vccd1
+ vccd1 _02240_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1299_X net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09668_ _02903_ _03629_ _04767_ _02940_ net442 vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__o32a_1
XANTENNA__07802__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ net1107 cpu.RF0.registers\[27\]\[3\] net881 vssd1 vssd1 vccd1 vccd1 _03910_
+ sky130_fd_sc_hd__and3_1
X_09599_ _04888_ _04889_ net277 vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ net2398 net138 net359 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13875__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__A1_N _03434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ net2118 net149 net367 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XANTENNA__07240__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13300_ clknet_leaf_30_clk cpu.RU0.next_FetchedData\[7\] net1208 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10512_ net1134 net1617 net914 _05643_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__a31o_1
XANTENNA__13105__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14280_ clknet_leaf_97_clk _01393_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11492_ net2597 net178 net376 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ clknet_leaf_44_clk _00411_ net1312 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10443_ net1130 net754 a1.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__or3b_2
XFILLER_0_61_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ clknet_leaf_52_clk net1643 net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ _01939_ _05477_ _05601_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__nor3_1
X_12113_ net744 _05987_ net557 vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__and3_4
XANTENNA__13255__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ clknet_leaf_51_clk _00273_ net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12145__B1 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14500__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12044_ cpu.LCD0.cnt_500hz\[0\] cpu.LCD0.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1 _05959_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09561__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09561__B2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net792 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13995_ clknet_leaf_86_clk _01108_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14650__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11933__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10459__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ clknet_leaf_20_clk _00135_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07712__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12877_ clknet_leaf_0_clk cpu.c0.next_count\[8\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14616_ clknet_leaf_52_clk net1530 net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09077__A0 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ net1951 net139 net334 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07088__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14547_ clknet_leaf_61_clk _01649_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_11759_ net1905 net148 net345 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__mux2_1
XANTENNA__08824__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478_ clknet_leaf_30_clk _00014_ net1207 vssd1 vssd1 vccd1 vccd1 cpu.RU0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08543__A _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14030__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ clknet_leaf_73_clk _00542_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11187__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08970_ cpu.RF0.registers\[9\]\[26\] net699 net650 cpu.RF0.registers\[14\]\[26\]
+ _04253_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__a221o_1
XANTENNA__14180__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07921_ net1030 cpu.RF0.registers\[22\]\[30\] net800 vssd1 vssd1 vccd1 vccd1 _03212_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10698__A0 cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__B _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12004__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ net1047 net634 net519 vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a21o_1
XANTENNA__06510__B cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ cpu.CU0.funct3\[1\] _01781_ cpu.CU0.bit30 cpu.CU0.funct3\[2\] vssd1 vssd1
+ vccd1 vccd1 _02094_ sky130_fd_sc_hd__or4bb_4
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
XFILLER_0_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07783_ cpu.RF0.registers\[15\]\[21\] net590 net565 cpu.RF0.registers\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a22o_1
XANTENNA__07325__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10032__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _04793_ _04794_ _04811_ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__o211a_2
XANTENNA__13898__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06734_ net1117 net1113 net1111 net1115 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07622__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _04687_ _04706_ net473 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06665_ a1.CPU_DAT_O\[1\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout252_A _05774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ cpu.RF0.registers\[18\]\[10\] net680 net666 _03693_ _03694_ vssd1 vssd1 vccd1
+ vccd1 _03695_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13128__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ net295 net298 _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09607__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06596_ cpu.LCD0.currentState\[5\] cpu.LCD0.nextState\[5\] _01965_ vssd1 vssd1 vccd1
+ vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ cpu.RF0.registers\[14\]\[12\] net650 _03624_ _03625_ net665 vssd1 vssd1 vccd1
+ vccd1 _03626_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12611__A1 cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09549__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07094__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ cpu.RF0.registers\[14\]\[15\] net649 net640 cpu.RF0.registers\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07217_ _02507_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ net940 cpu.RF0.registers\[2\]\[21\] net855 vssd1 vssd1 vccd1 vccd1 _03488_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14523__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07069__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08043__A1 cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ cpu.RF0.registers\[0\]\[11\] net620 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08594__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__Y _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ cpu.RF0.registers\[21\]\[18\] net593 net588 cpu.RF0.registers\[1\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1007 net1011 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_4
X_10090_ _05360_ _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__and2_1
Xfanout1018 cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
Xfanout1029 net1033 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677__1399 vssd1 vssd1 vccd1 vccd1 _14677__1399/HI net1399 sky130_fd_sc_hd__conb_1
XFILLER_0_92_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__C net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ net2676 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13780_ clknet_leaf_70_clk _00893_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ _03041_ net533 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nor2_1
XANTENNA__07306__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ cpu.f0.state\[7\] net497 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12662_ net2280 net2186 net1009 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14053__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14401_ clknet_leaf_17_clk _01512_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_11613_ net1736 net199 net358 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XANTENNA__12602__A1 cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__Q cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _05155_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ clknet_leaf_56_clk _01445_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07085__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net1921 net215 net367 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14263_ clknet_leaf_65_clk _01376_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ net2061 net225 net377 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ clknet_leaf_63_clk _00394_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ cpu.f0.i\[25\] net268 vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14194_ clknet_leaf_60_clk _01307_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09782__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11928__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ clknet_leaf_48_clk _00325_ net1355 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[109\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10832__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ _05589_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nand2_1
XANTENNA__07707__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ clknet_leaf_50_clk net2227 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10288_ cpu.f0.i\[17\] net541 _05526_ net526 vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a31o_1
XANTENNA__08337__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ net2874 net128 net310 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__mux2_1
XANTENNA__10144__A2 _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11663__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ clknet_leaf_93_clk _01091_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07442__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12929_ clknet_leaf_28_clk _00118_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10852__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06450_ net2671 _01826_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[6\] sky130_fd_sc_hd__xor2_1
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06381_ cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13420__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14546__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ net935 cpu.RF0.registers\[8\]\[23\] net870 vssd1 vssd1 vccd1 vccd1 _03411_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08273__A1 cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08051_ net939 cpu.RF0.registers\[14\]\[25\] net838 vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06505__B cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ net955 cpu.RF0.registers\[15\]\[23\] net825 vssd1 vssd1 vccd1 vccd1 _02293_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_71_clk_X clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13570__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload37_A clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__X _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12109__B1 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08328__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07904_ net523 _03192_ _03194_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_leaf_86_clk_X clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ net937 cpu.RF0.registers\[14\]\[17\] net837 vssd1 vssd1 vccd1 vccd1 _04175_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10043__A cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10135__A2 _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__X _04682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07835_ cpu.RF0.registers\[22\]\[24\] net604 net570 cpu.RF0.registers\[10\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__a22o_1
XANTENNA__10978__A _02981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07766_ net962 cpu.RF0.registers\[11\]\[21\] net776 vssd1 vssd1 vccd1 vccd1 _03057_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14076__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _03594_ _03629_ net468 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__mux2_1
XANTENNA__06894__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ net1113 net1110 net1116 net1114 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__and4b_2
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ net1031 cpu.RF0.registers\[29\]\[17\] net791 vssd1 vssd1 vccd1 vccd1 _02988_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07303__A3 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08500__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09436_ _03019_ _04402_ _04725_ net298 net291 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06648_ net2270 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[16\] sky130_fd_sc_hd__and2_1
XFILLER_0_52_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_clk_X clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout801_A _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ _04525_ _04530_ net475 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ cpu.LCD0.cnt_500hz\[0\] cpu.LCD0.cnt_500hz\[1\] cpu.LCD0.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__nand3_1
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08318_ net1089 cpu.RF0.registers\[17\]\[12\] net883 vssd1 vssd1 vccd1 vccd1 _03609_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08183__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_50 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ net305 _04583_ _04586_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10071__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13913__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _03538_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1331_X net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ net2175 net179 net405 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11020__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _05458_ _05462_ _05471_ net132 net715 vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ net1744 net168 net411 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ net718 net135 _05408_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a22o_1
X_10073_ cpu.IM0.address_IM\[20\] _03042_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xor2_1
XANTENNA__07527__B1 _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ clknet_leaf_102_clk _01014_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13037__Q cpu.LCD0.row_1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_84_clk _00945_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07262__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ clknet_leaf_75_clk _00876_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10975_ _02433_ _05849_ _05851_ net532 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__o211a_2
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13443__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12714_ cpu.LCD0.row_2\[116\] cpu.LCD0.row_2\[108\] net1008 vssd1 vssd1 vccd1 vccd1
+ _01707_ sky130_fd_sc_hd__mux2_1
XANTENNA__14569__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ clknet_leaf_85_clk _00807_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ net2214 net2448 net1007 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07058__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ cpu.DM0.data_i\[4\] _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13593__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire240 _04753_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
X_14315_ clknet_leaf_86_clk _01428_ net1272 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08524__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__A2 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ net1949 net158 net370 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__mux2_1
XANTENNA__13981__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 cpu.RF0.registers\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ clknet_leaf_5_clk _01359_ net1148 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ net2591 net153 net378 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11658__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ net1125 _05622_ net264 net1999 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14177_ clknet_leaf_60_clk _01290_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11389_ net2645 net182 net387 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13128_ clknet_leaf_49_clk _00308_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_13059_ clknet_leaf_53_clk net2179 net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 cpu.RF0.registers\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1360 net1362 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__clkbuf_4
Xfanout1371 net1385 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__clkbuf_2
Xfanout1382 net1383 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11393__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ net964 cpu.RF0.registers\[5\]\[13\] net796 vssd1 vssd1 vccd1 vccd1 _02911_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_50_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ net1052 cpu.RF0.registers\[20\]\[8\] net783 vssd1 vssd1 vccd1 vccd1 _02842_
+ sky130_fd_sc_hd__and3_1
X_06502_ cpu.K0.keyvalid cpu.f0.state\[5\] _01890_ vssd1 vssd1 vccd1 vccd1 _01892_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07297__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ net980 cpu.RF0.registers\[9\]\[5\] net760 vssd1 vssd1 vccd1 vccd1 _02773_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12290__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09221_ net449 _04511_ _04510_ _04384_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o211ai_1
X_06433_ cpu.c0.count\[11\] cpu.c0.count\[12\] _01840_ vssd1 vssd1 vccd1 vccd1 _01843_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13936__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12518__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ net480 _04371_ _04377_ _04382_ _04390_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09099__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06364_ cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14676__1398 vssd1 vssd1 vccd1 vccd1 _14676__1398/HI net1398 sky130_fd_sc_hd__conb_1
XFILLER_0_72_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08103_ cpu.RF0.registers\[8\]\[22\] net708 _03376_ _03377_ _03379_ vssd1 vssd1 vccd1
+ vccd1 _03394_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09994__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09083_ net464 net449 net437 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_20_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10038__A cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__B_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ cpu.RF0.registers\[23\]\[24\] net671 _03310_ _03311_ _03312_ vssd1 vssd1
+ vccd1 vccd1 _03325_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09827__A _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold810 cpu.LCD0.row_1\[50\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06803__X _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold821 _00256_ vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 cpu.LCD0.row_2\[118\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11568__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold843 cpu.RF0.registers\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__B _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 cpu.RF0.registers\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 cpu.RF0.registers\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 cpu.RF0.registers\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06889__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold887 cpu.RF0.registers\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 _00251_ vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13316__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net629 _04813_ net931 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout584_A _02173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08936_ net938 cpu.RF0.registers\[13\]\[27\] net849 vssd1 vssd1 vccd1 vccd1 _04227_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12540__X _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1510 cpu.f0.num\[30\] vssd1 vssd1 vccd1 vccd1 net2916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06980__B2 cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1521 cpu.RF0.registers\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net2927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1532 cpu.LCD0.row_2\[11\] vssd1 vssd1 vccd1 vccd1 net2938 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ cpu.IM0.address_IM\[16\] net551 _04156_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout751_A _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13466__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A _02041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__Y _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ cpu.RF0.registers\[11\]\[22\] net567 _03082_ _03090_ _03096_ vssd1 vssd1
+ vccd1 vccd1 _03109_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_93_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08798_ _04088_ net441 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ _03025_ _03026_ _03038_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07513__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ _05688_ _05717_ _05718_ net1017 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1
+ vccd1 _05719_ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12281__A2 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09419_ net450 _04471_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__or2_2
XANTENNA__07810__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ net2727 cpu.LCD0.row_1\[105\] net906 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12430_ cpu.DM0.data_i\[23\] net535 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09985__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net1122 net1526 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13320__Q cpu.DM0.data_i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ clknet_leaf_73_clk _01213_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13392__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ net2000 net218 net394 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__mux2_1
XANTENNA__06713__X _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ _06105_ _06157_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__nor2_1
XANTENNA__07460__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14031_ clknet_leaf_81_clk _01144_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11478__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ net2719 net226 net405 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10989__B1_N net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07257__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11174_ net2797 net241 net412 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__mux2_1
XANTENNA__14241__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__A2_N net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _05346_ _05362_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__nand3_1
XANTENNA__13809__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07691__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _02004_ _05146_ _05329_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08712__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14391__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08088__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08519__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13959__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ clknet_leaf_64_clk _00928_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11941__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13746_ clknet_leaf_70_clk _00859_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07279__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ net273 _05855_ _05856_ net925 net1662 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12272__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13677_ clknet_leaf_101_clk _00790_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ _05321_ _05811_ net719 vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__mux2_1
XANTENNA__12983__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ net2622 net2497 net1006 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10035__A1 cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ _06322_ _06323_ _06324_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__or4_4
XANTENNA__09976__B2 _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13339__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold106 cpu.DM0.readdata\[15\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 net99 vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 cpu.LCD0.row_2\[122\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11388__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 cpu.f0.write_data\[23\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ clknet_leaf_73_clk _01342_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07739__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout608 _02141_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_8
XFILLER_0_10_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13489__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _04034_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08951__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ net544 _02272_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14268__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ cpu.RF0.registers\[28\]\[0\] net1096 net868 vssd1 vssd1 vccd1 vccd1 _04012_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10256__C_N net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12012__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ net1102 cpu.RF0.registers\[26\]\[2\] _02025_ vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10510__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07603_ _02890_ _02891_ _02892_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__or4_1
X_08583_ net1100 cpu.RF0.registers\[24\]\[4\] net871 vssd1 vssd1 vccd1 vccd1 _03874_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07333__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07534_ _02821_ _02822_ _02823_ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__or4_1
XANTENNA__12263__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07630__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07465_ net523 _02754_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout332_A _05938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14114__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09204_ _04413_ _04488_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__nor2_1
X_06416_ cpu.c0.count\[16\] _01824_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07690__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ net971 cpu.RF0.registers\[6\]\[0\] net803 vssd1 vssd1 vccd1 vccd1 _02687_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08164__C net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09135_ _04422_ _04425_ net455 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13140__Q cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1241_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1339_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09557__A _02865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09066_ cpu.RF0.registers\[0\]\[31\] net617 _04351_ _04356_ vssd1 vssd1 vccd1 vccd1
+ _04357_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_92_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08461__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14264__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09719__A1 _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ net1099 cpu.RF0.registers\[27\]\[24\] net879 vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout799_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 cpu.RF0.registers\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 cpu.RF0.registers\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold662 cpu.RF0.registers\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07077__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 cpu.RF0.registers\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 cpu.RF0.registers\[4\]\[11\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold695 cpu.RF0.registers\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07508__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _05247_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nand2_2
XANTENNA__10930__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11012__B1_N net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _04128_ _04198_ _04207_ _04209_ _04126_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__o311a_1
XANTENNA__07805__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ _05173_ _05174_ _05171_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a21o_1
Xhold1340 cpu.RF0.registers\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08155__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11930_ net2207 net237 net320 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
Xhold1351 cpu.RF0.registers\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 cpu.f0.data_adr\[26\] vssd1 vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1384 cpu.RF0.registers\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 cpu.K0.code\[0\] vssd1 vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11861_ net1877 net137 net330 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11027__B1_N net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ clknet_leaf_9_clk _00713_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10812_ cpu.IM0.address_IM\[28\] net1014 net285 _05755_ vssd1 vssd1 vccd1 vccd1 _05756_
+ sky130_fd_sc_hd__a22o_1
X_14580_ clknet_leaf_46_clk net2341 net1356 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12254__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net1598 net148 net338 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13531_ clknet_leaf_12_clk _00644_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10743_ net1604 net559 net537 _05706_ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13462_ clknet_leaf_59_clk _00575_ net1348 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09407__A0 _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net2720 net2679 net910 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XANTENNA__07681__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10017__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12413_ cpu.CU0.funct3\[0\] cpu.DM0.data_i\[15\] _01848_ _02095_ _06222_ vssd1 vssd1
+ vccd1 vccd1 _06230_ sky130_fd_sc_hd__a41o_1
X_13393_ clknet_leaf_79_clk _00506_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12344_ net2841 _06212_ net1368 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_75_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08802__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12275_ _06152_ _06154_ _06156_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13631__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ clknet_leaf_86_clk _01127_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11226_ net2792 _05827_ net406 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
XANTENNA__07418__C net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net2184 net183 net416 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10840__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ net126 _05378_ _05375_ net627 vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_88_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13781__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ net1661 net187 net423 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
X_14675__1397 vssd1 vssd1 vccd1 vccd1 _14675__1397/HI net1397 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10039_ _05312_ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07153__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13011__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14137__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12245__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06992__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ clknet_leaf_63_clk _00842_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07250_ cpu.RF0.registers\[14\]\[9\] net576 _02518_ _02522_ _02526_ vssd1 vssd1 vccd1
+ vccd1 _02541_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13161__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14287__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10008__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09949__A1 cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07181_ _02438_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08281__A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09096__B _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10316__A cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06513__B cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14449__RESET_B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout405 _05919_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_4
XANTENNA__07328__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_6
X_09822_ _04475_ _04677_ _04929_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__o22ai_1
XANTENNA__11846__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout427 _05911_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_4
Xfanout438 _04323_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_4
Xfanout449 net452 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
XANTENNA__07625__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ net481 _04835_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__nor2_1
X_06965_ cpu.RF0.registers\[29\]\[25\] net601 _02252_ _02255_ vssd1 vssd1 vccd1 vccd1
+ _02256_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout282_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _03992_ _03993_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand3_1
X_09684_ net476 _03964_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__or2_1
X_06896_ net971 net759 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ cpu.RF0.registers\[11\]\[3\] net688 _02033_ cpu.RF0.registers\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07063__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1191_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11581__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1289_A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ cpu.RF0.registers\[5\]\[5\] net704 net649 cpu.RF0.registers\[14\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13504__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ net981 cpu.RF0.registers\[8\]\[6\] net814 vssd1 vssd1 vccd1 vccd1 _02808_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _03784_ _03785_ _03786_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07448_ net1056 cpu.RF0.registers\[21\]\[1\] net797 vssd1 vssd1 vccd1 vccd1 _02739_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_94_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07379_ cpu.RF0.registers\[5\]\[2\] net602 _02658_ _02659_ _02666_ vssd1 vssd1 vccd1
+ vccd1 _02670_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10925__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1244_X net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ _04379_ _04391_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or2_4
X_10390_ net1021 net268 vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__nand2_1
XANTENNA__07415__A2 _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08622__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ net952 cpu.RF0.registers\[9\]\[31\] net756 vssd1 vssd1 vccd1 vccd1 _04340_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12966__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10970__A2 _05863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ cpu.LCD0.cnt_500hz\[7\] _05966_ cpu.LCD0.cnt_500hz\[8\] vssd1 vssd1 vccd1
+ vccd1 _05968_ sky130_fd_sc_hd__a21o_1
Xhold470 cpu.RF0.registers\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold481 cpu.RF0.registers\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07238__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ net1729 net928 net276 _05893_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a22o_1
Xhold492 _01702_ vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14119__RESET_B net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07094__X _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net951 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_2
Xfanout961 net984 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_2
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_1
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_2
Xfanout994 net996 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13034__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ clknet_leaf_28_clk _00151_ net1183 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1170 cpu.RF0.registers\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net2189 net207 net322 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
Xhold1181 cpu.RF0.registers\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1192 cpu.RF0.registers\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ clknet_leaf_33_clk _00024_ net1245 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12587__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14632_ clknet_leaf_31_clk _01733_ net1202 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_11844_ net1976 net198 net330 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
XANTENNA__12227__A2 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14563_ clknet_leaf_61_clk net2635 net1345 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07701__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ net2245 net212 net339 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10789__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08300__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10726_ a1.ADR_I\[3\] net559 net537 _05694_ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__a22o_1
X_13514_ clknet_leaf_100_clk _00627_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ clknet_leaf_34_clk _01596_ net1251 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[5\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13445_ clknet_leaf_9_clk _00558_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10835__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ net2111 cpu.LCD0.row_1\[71\] net903 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload15 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_58_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload26 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload26/X sky130_fd_sc_hd__clkbuf_4
X_13376_ clknet_leaf_8_clk _00489_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload37 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload37/X sky130_fd_sc_hd__clkbuf_4
X_10588_ _05682_ cpu.LCD0.row_1\[5\] net896 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
XANTENNA__09800__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload48 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload59 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12327_ cpu.LCD0.cnt_20ms\[8\] _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12258_ cpu.LCD0.row_2\[102\] _06018_ _06033_ cpu.LCD0.row_2\[78\] vssd1 vssd1 vccd1
+ vccd1 _06153_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11666__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ net2386 net228 net409 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
X_12189_ cpu.LCD0.row_2\[107\] _06012_ _06030_ cpu.LCD0.row_1\[43\] _06086_ vssd1
+ vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07445__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06987__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ net1115 net1117 net1111 net1113 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__and4b_2
XFILLER_0_56_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13527__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06681_ a1.CPU_DAT_O\[17\] net889 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[17\]
+ sky130_fd_sc_hd__and2_1
X_08420_ net1079 cpu.RF0.registers\[22\]\[9\] net851 vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12218__A2 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ net940 cpu.RF0.registers\[3\]\[11\] net835 vssd1 vssd1 vccd1 vccd1 _03642_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09095__A1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06508__B cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13677__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07302_ cpu.RF0.registers\[22\]\[4\] net604 net583 cpu.RF0.registers\[6\]\[4\] _02592_
+ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a221o_1
X_08282_ net1082 cpu.RF0.registers\[26\]\[13\] net860 vssd1 vssd1 vccd1 vccd1 _03573_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07645__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload67_A clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinv_8
X_07233_ net955 cpu.RF0.registers\[13\]\[9\] net790 vssd1 vssd1 vccd1 vccd1 _02524_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12085__X _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07179__X _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07164_ net1043 cpu.RF0.registers\[26\]\[11\] net787 vssd1 vssd1 vccd1 vccd1 _02455_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08070__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07095_ cpu.RF0.registers\[23\]\[14\] net613 net586 cpu.RF0.registers\[4\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1037_A cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout213 net215 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
Xfanout224 _05786_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
Xfanout235 _05781_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xfanout246 _05776_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_1
XANTENNA__06897__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _06264_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
X_09805_ net493 _04552_ _05087_ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a31o_2
Xfanout268 net271 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
X_07997_ cpu.RF0.registers\[29\]\[28\] net672 net646 cpu.RF0.registers\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net482 net436 _04973_ _04397_ net290 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__o221a_1
X_06948_ cpu.RF0.registers\[1\]\[26\] net588 _02214_ _02221_ _02223_ vssd1 vssd1 vccd1
+ vccd1 _02239_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09322__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _02410_ _03534_ _04946_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or3b_1
XANTENNA__14452__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10468__B2 a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ net962 cpu.RF0.registers\[1\]\[27\] net805 vssd1 vssd1 vccd1 vccd1 _02170_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ net1107 cpu.RF0.registers\[23\]\[3\] net845 vssd1 vssd1 vccd1 vccd1 _03909_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ _04384_ _04823_ _04885_ net486 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a22o_1
XANTENNA__07884__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08617__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ net1105 cpu.RF0.registers\[27\]\[5\] net881 vssd1 vssd1 vccd1 vccd1 _03840_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07521__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12090__B1 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net2475 net156 net366 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
X_10511_ net40 net919 vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11491_ cpu.RF0.registers\[14\]\[23\] net153 net374 vssd1 vssd1 vccd1 vccd1 _00911_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13230_ clknet_leaf_44_clk _00410_ net1312 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14674__1396 vssd1 vssd1 vccd1 vccd1 _14674__1396/HI net1396 sky130_fd_sc_hd__conb_1
X_10442_ net1130 a1.prev_BUSY_O net752 vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__and3b_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08352__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08597__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ clknet_leaf_48_clk _00341_ net1355 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[125\]
+ sky130_fd_sc_hd__dfstp_1
X_10373_ _01861_ _01864_ _05603_ net1130 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12112_ cpu.LCD0.row_2\[48\] _06011_ _06012_ cpu.LCD0.row_2\[104\] _06010_ vssd1
+ vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a221o_1
X_13092_ clknet_leaf_50_clk _00272_ net1382 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ cpu.LCD0.cnt_500hz\[0\] net502 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__and2b_1
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_4
Xfanout791 net792 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06780__C1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ clknet_leaf_101_clk _01107_ net1213 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09313__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__B2 a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12945_ clknet_leaf_20_clk _00134_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12876_ clknet_leaf_0_clk cpu.c0.next_count\[7\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07875__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ clknet_leaf_55_clk net1432 net1367 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11827_ net2494 net140 net336 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__mux2_1
XANTENNA__07431__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__A1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14546_ clknet_leaf_51_clk _01648_ net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_11758_ net2592 net155 net342 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ cpu.LCD0.row_1\[115\] net1600 net897 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14477_ clknet_leaf_33_clk _01587_ net1250 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09639__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11689_ net2849 net154 net350 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13428_ clknet_leaf_70_clk _00541_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12384__B2 cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ clknet_leaf_82_clk _00472_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07727__X _03018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11396__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ net957 cpu.RF0.registers\[10\]\[30\] net787 vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10147__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07851_ cpu.RF0.registers\[0\]\[24\] net618 _03135_ _03141_ vssd1 vssd1 vccd1 vccd1
+ _03142_ sky130_fd_sc_hd__o22a_4
XANTENNA__14475__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__A_N net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ cpu.CU0.funct3\[1\] _01781_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__or2_1
XANTENNA__12917__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ _03069_ _03070_ _03071_ _03072_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__or4_1
X_09521_ net278 _04713_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__nand2_1
XANTENNA__07462__X _02753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06733_ net1087 net883 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__and2_2
XANTENNA__07903__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07315__A1 cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07315__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ net306 _04742_ _04697_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__o21a_1
X_06664_ a1.CPU_DAT_O\[0\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12020__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07866__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ cpu.RF0.registers\[1\]\[10\] net714 _03670_ _03677_ _03686_ vssd1 vssd1 vccd1
+ vccd1 _03694_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09383_ _02348_ _04123_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nand2_1
X_06595_ _01756_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout245_A _05776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ cpu.RF0.registers\[4\]\[12\] net677 _03602_ _03606_ _03612_ vssd1 vssd1 vccd1
+ vccd1 _03625_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07079__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ cpu.RF0.registers\[30\]\[15\] net660 net647 cpu.RF0.registers\[21\]\[15\]
+ _03543_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__a221o_1
XANTENNA__09549__B _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08291__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout412_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1154_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ _02474_ _02506_ net544 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ net939 cpu.RF0.registers\[8\]\[21\] net870 vssd1 vssd1 vccd1 vccd1 _03487_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12375__B2 cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12690__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ _01851_ _02123_ cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1321_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ cpu.RF0.registers\[16\]\[18\] net581 _02352_ _02356_ _02365_ vssd1 vssd1
+ vccd1 vccd1 _02369_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout781_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 net1011 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_2
Xfanout1019 cpu.f0.i\[22\] vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07516__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13842__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _04397_ _04393_ _04970_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__mux2_1
X_10991_ a1.CPU_DAT_I\[19\] net929 _05846_ _05879_ vssd1 vssd1 vccd1 vccd1 _00427_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08503__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ net528 _01942_ _01760_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_2_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08347__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ cpu.LCD0.row_2\[63\] net2109 net1007 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__mux2_1
XANTENNA__13992__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11612_ net2084 net210 net358 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
X_14400_ clknet_leaf_21_clk _01511_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ cpu.IM0.address_IM\[0\] _02682_ _05153_ _05154_ vssd1 vssd1 vccd1 vccd1 _06351_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08644__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__X _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ net2059 net218 net366 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
X_14331_ clknet_leaf_56_clk _01444_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10238__X _05490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13222__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14348__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14262_ clknet_leaf_59_clk _01375_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ net2373 net230 net377 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XANTENNA__07490__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13213_ clknet_leaf_8_clk _00393_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14134__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10425_ _01816_ net269 _05630_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12366__B2 cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09231__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ clknet_leaf_77_clk _01306_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13144_ clknet_leaf_48_clk _00324_ net1362 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[108\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ cpu.f0.i\[27\] _05585_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14498__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13075_ clknet_leaf_51_clk net2053 net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ net1998 _05531_ net727 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12026_ net2584 net137 net310 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__mux2_1
XANTENNA__11944__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09298__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ clknet_leaf_14_clk _01090_ net1240 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ clknet_leaf_26_clk _00117_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10301__B1 _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07161__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ clknet_leaf_23_clk _00078_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_06380_ cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08554__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14529_ clknet_leaf_49_clk _01631_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08273__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ net1087 cpu.RF0.registers\[23\]\[25\] net847 vssd1 vssd1 vccd1 vccd1 _03341_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10308__B cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13715__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07001_ net955 cpu.RF0.registers\[3\]\[23\] net820 vssd1 vssd1 vccd1 vccd1 _02292_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09222__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06802__A cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12109__B2 cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08981__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08720__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ cpu.IM0.address_IM\[27\] net552 _04241_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_
+ sky130_fd_sc_hd__a22o_4
XANTENNA__13865__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06521__B cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ net544 _03193_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or2_1
X_08883_ net935 cpu.RF0.registers\[12\]\[17\] net867 vssd1 vssd1 vccd1 vccd1 _04174_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07336__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ cpu.RF0.registers\[29\]\[24\] net601 net596 cpu.RF0.registers\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10978__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07633__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14673__1395 vssd1 vssd1 vccd1 vccd1 _14673__1395/HI net1395 sky130_fd_sc_hd__conb_1
X_07765_ net962 cpu.RF0.registers\[6\]\[21\] net801 vssd1 vssd1 vccd1 vccd1 _03056_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout362_A _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ _03534_ _03564_ net464 vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__mux2_1
X_06716_ net946 net884 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__and2_4
XANTENNA__12293__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07839__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ net1027 cpu.RF0.registers\[21\]\[17\] net795 vssd1 vssd1 vccd1 vccd1 _02987_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ net293 _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor2_1
XANTENNA__08167__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07071__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06647_ a1.CPU_DAT_O\[15\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[15\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__13245__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09366_ _04413_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__or2_1
X_06578_ cpu.LCD0.cnt_500hz\[0\] cpu.LCD0.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1 _01953_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08464__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ net1086 cpu.RF0.registers\[22\]\[12\] net851 vssd1 vssd1 vccd1 vccd1 _03608_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_40 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ net296 _04587_ _04585_ _04584_ _04562_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_51 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _03534_ _03537_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10071__A2 _04683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13395__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14640__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ cpu.RF0.registers\[0\]\[20\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03470_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__10359__B1 _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _05458_ _05462_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a21o_1
XANTENNA__07808__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net2292 net184 net412 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08972__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _05405_ _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10234__A cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A2_N _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ _05344_ _05345_ cpu.IM0.address_IM\[19\] net1023 vssd1 vssd1 vccd1 vccd1
+ _00042_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13318__Q cpu.DM0.data_i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ clknet_leaf_88_clk _01013_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07543__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ clknet_leaf_79_clk _00944_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14020__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11087__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ _02433_ net516 vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__and2b_1
X_13762_ clknet_leaf_10_clk _00875_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12713_ net2262 net2149 net1002 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13693_ clknet_leaf_88_clk _00806_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14170__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12644_ net2233 cpu.LCD0.row_2\[38\] net1005 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13738__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10598__A0 cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12575_ cpu.DM0.data_i\[6\] cpu.DM0.data_i\[0\] cpu.DM0.data_i\[1\] _06338_ vssd1
+ vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09452__A1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08255__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11004__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14314_ clknet_leaf_102_clk _01427_ net1215 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11526_ net2040 net161 net372 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11939__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ net1919 net165 net378 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
X_14245_ clknet_leaf_9_clk _01358_ net1166 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10843__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__X _06082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13888__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ cpu.f0.i\[16\] net268 vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nand2_1
X_14176_ clknet_leaf_9_clk _01289_ net1162 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11388_ net2001 net170 net386 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__mux2_1
X_13127_ clknet_leaf_46_clk net1820 net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_10339_ net2768 net724 _05575_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_81_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13118__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ clknet_leaf_52_clk net2337 net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07156__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1364 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__clkbuf_2
X_12009_ net2087 net199 net311 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__mux2_1
Xfanout1361 net1362 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1372 net1377 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__clkbuf_4
Xfanout1383 net1384 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06995__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13268__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ net1052 cpu.RF0.registers\[28\]\[8\] net767 vssd1 vssd1 vccd1 vccd1 _02841_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14513__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06501_ cpu.K0.keyvalid _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ net1060 cpu.RF0.registers\[25\]\[5\] net760 vssd1 vssd1 vccd1 vccd1 _02772_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09691__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09691__B2 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _03372_ _04276_ net465 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06432_ cpu.c0.count\[13\] cpu.c0.count\[12\] cpu.c0.count\[14\] _01841_ vssd1 vssd1
+ vccd1 vccd1 _01842_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08284__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12578__A1 cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__B cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14056__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ _04427_ _04441_ net486 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
X_06363_ cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__inv_2
XANTENNA__10589__A0 cpu.f0.write_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ cpu.RF0.registers\[29\]\[22\] net672 _03382_ _03383_ _03385_ vssd1 vssd1
+ vccd1 vccd1 _03393_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09082_ net465 net448 _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ cpu.RF0.registers\[14\]\[24\] net649 _03309_ _03315_ _03319_ vssd1 vssd1
+ vccd1 vccd1 _03324_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11849__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12093__X _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__B _05086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold800 cpu.RF0.registers\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 _00274_ vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout208_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 cpu.RF0.registers\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _01709_ vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__B2 a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold844 cpu.RF0.registers\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 cpu.f0.num\[26\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold866 cpu.RF0.registers\[4\]\[6\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12750__B2 cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 cpu.LCD0.row_1\[42\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold888 cpu.RF0.registers\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net125 _05262_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a21o_1
Xhold899 cpu.RF0.registers\[8\]\[17\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10761__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ net1083 cpu.RF0.registers\[22\]\[27\] net851 vssd1 vssd1 vccd1 vccd1 _04226_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14043__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 cpu.f0.num\[24\] vssd1 vssd1 vccd1 vccd1 net2906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout577_A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1511 cpu.RF0.registers\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net2917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 net124 vssd1 vssd1 vccd1 vccd1 net2928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 a1.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net2939 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ cpu.RF0.registers\[0\]\[16\] net661 net547 vssd1 vssd1 vccd1 vccd1 _04157_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08182__A1 _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08459__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07817_ cpu.RF0.registers\[24\]\[22\] net608 _03085_ _03088_ _03089_ vssd1 vssd1
+ vccd1 vccd1 _03108_ sky130_fd_sc_hd__a2111o_1
X_08797_ _02383_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14193__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12266__B1 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ cpu.RF0.registers\[20\]\[20\] _02160_ net581 cpu.RF0.registers\[16\]\[20\]
+ _03028_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout911_A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ net953 cpu.RF0.registers\[5\]\[16\] net795 vssd1 vssd1 vccd1 vccd1 _02970_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10928__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _04466_ _04473_ net450 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__mux2_1
X_10690_ net2739 cpu.LCD0.row_1\[104\] net910 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XANTENNA__07693__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08237__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ _04578_ _04618_ _04638_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a21o_2
XANTENNA__10229__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12360_ net1122 net1954 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__and2_1
XANTENNA__09985__A2 _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08922__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ net1653 net221 net396 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ cpu.LCD0.row_2\[63\] _06000_ _06009_ cpu.LCD0.row_1\[111\] _06184_ vssd1
+ vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09198__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14030_ clknet_leaf_1_clk _01143_ net1139 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11242_ net2552 net230 net405 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__mux2_1
XANTENNA__12741__A1 cpu.f0.write_data\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11173_ net2889 net246 net412 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07212__A3 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ _05371_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__and3_1
XANTENNA__06971__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13410__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _05326_ _05328_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__nand2_1
XANTENNA__14536__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07273__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ clknet_leaf_70_clk _00927_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12257__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_70_clk_X clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13560__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ clknet_leaf_76_clk _00858_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10838__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ net985 cpu.f0.write_data\[9\] vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11480__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ clknet_leaf_80_clk _00789_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ cpu.DM0.readdata\[17\] _04734_ net734 vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ cpu.LCD0.row_2\[29\] cpu.LCD0.row_2\[21\] net1000 vssd1 vssd1 vccd1 vccd1
+ _01620_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08228__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ _01870_ _01890_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06904__X _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11509_ net1735 net220 net372 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__mux2_1
XANTENNA__09647__B _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold107 a1.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
X_14672__1394 vssd1 vssd1 vccd1 vccd1 _14672__1394/HI net1394 sky130_fd_sc_hd__conb_1
X_12489_ _05506_ net257 cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold118 _00156_ vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10991__B1 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__B1 _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold129 _01713_ vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ clknet_leaf_70_clk _01341_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159_ clknet_leaf_87_clk _01272_ net1287 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout609 _02139_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_8
XANTENNA__08400__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ cpu.IG0.Instr\[25\] net633 net519 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_23_clk_X clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13090__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09382__B _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ cpu.RF0.registers\[8\]\[0\] net946 net871 vssd1 vssd1 vccd1 vccd1 _04011_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08279__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__A cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1191 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_2
Xfanout1191 net1211 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_2
X_08651_ cpu.RF0.registers\[4\]\[2\] net679 _03939_ _03940_ _03941_ vssd1 vssd1 vccd1
+ vccd1 _03942_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07614__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07602_ cpu.RF0.registers\[13\]\[12\] net597 net593 cpu.RF0.registers\[21\]\[12\]
+ _02871_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a221o_1
XANTENNA__12248__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08582_ cpu.RF0.registers\[7\]\[4\] net652 net647 cpu.RF0.registers\[21\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a22o_1
XANTENNA__09113__B1 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14237__RESET_B net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ cpu.RF0.registers\[10\]\[6\] net570 _02800_ _02803_ _02809_ vssd1 vssd1 vccd1
+ vccd1 _02824_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload97_A clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08467__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12529__A cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout158_A _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ net525 _02719_ _02720_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__nand3_4
XFILLER_0_91_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06415_ cpu.c0.count\[6\] _01826_ cpu.c0.count\[7\] vssd1 vssd1 vccd1 vccd1 _01828_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09203_ net495 _03234_ _04492_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07395_ cpu.RF0.registers\[24\]\[0\] net607 _02683_ _02684_ _02685_ vssd1 vssd1 vccd1
+ vccd1 _02686_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10049__A cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _04423_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__B1 _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14409__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11579__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09065_ _04352_ _04353_ _04354_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or4_1
XANTENNA__09557__B _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13872__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ net947 cpu.RF0.registers\[6\]\[24\] net852 vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold630 cpu.RF0.registers\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 cpu.RF0.registers\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 cpu.RF0.registers\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold663 cpu.RF0.registers\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10734__A0 cpu.f0.data_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold674 cpu.RF0.registers\[16\]\[6\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13433__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 cpu.RF0.registers\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold696 cpu.RF0.registers\[6\]\[30\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout861_A _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net440 _04125_ _04089_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o21ai_1
X_09898_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__or2_1
XANTENNA__08189__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1330 cpu.RF0.registers\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 cpu.RF0.registers\[14\]\[5\] vssd1 vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13583__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1352 cpu.RF0.registers\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09711__D_N _05001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ cpu.RF0.registers\[13\]\[16\] net659 _04137_ _04138_ _04139_ vssd1 vssd1
+ vccd1 vccd1 _04140_ sky130_fd_sc_hd__a2111o_1
Xhold1363 cpu.RF0.registers\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07524__C net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__A1 cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1374 cpu.RF0.registers\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 cpu.RF0.registers\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12239__B1 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1396 cpu.RF0.registers\[13\]\[10\] vssd1 vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
X_11860_ net2780 net141 net333 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10811_ cpu.f0.data_adr\[28\] _04716_ net993 vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__mux2_1
X_11791_ net1761 net157 net338 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ clknet_leaf_93_clk _00643_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ cpu.IM0.address_IM\[8\] net1014 net286 _05705_ vssd1 vssd1 vccd1 vccd1 _05706_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08355__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10673_ cpu.LCD0.row_1\[79\] net2644 net902 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13461_ clknet_leaf_73_clk _00574_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09407__A1 _03300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12412_ net1614 net732 _06229_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__o21a_1
XANTENNA__10017__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14089__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ clknet_leaf_75_clk _00505_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11489__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12343_ cpu.LCD0.cnt_20ms\[14\] _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10973__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08630__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12274_ cpu.LCD0.row_1\[126\] _06014_ _06159_ _06168_ _01961_ vssd1 vssd1 vccd1 vccd1
+ _06169_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08090__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ net1975 net163 net406 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__mux2_1
X_14013_ clknet_leaf_68_clk _01126_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12190__A2 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net1811 net171 net414 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
XANTENNA__06900__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13926__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10107_ _05376_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ net2927 net192 net422 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10038_ cpu.IM0.address_IM\[17\] _02984_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__A1 cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08697__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11952__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12950__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ net2395 net157 net314 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__mux2_1
X_13728_ clknet_leaf_3_clk _00841_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13306__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07121__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ clknet_leaf_13_clk _00772_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09949__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ cpu.CU0.opcode\[6\] cpu.IG0.Instr\[7\] _01850_ _02004_ cpu.IG0.Instr\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11399__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13456__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10964__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09945__X _05229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout406 _05918_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
X_09821_ _02383_ net434 net288 _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__o211a_1
Xfanout417 _05916_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09393__A _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 _05911_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_6
Xfanout439 _04194_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload12_A clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _05032_ _05039_ _05042_ _05035_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__or4b_4
XANTENNA__12023__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06964_ cpu.RF0.registers\[28\]\[25\] net577 _02253_ _02254_ vssd1 vssd1 vccd1 vccd1
+ _02255_ sky130_fd_sc_hd__a211o_1
X_08703_ _02122_ net462 net456 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a21o_1
X_09683_ net482 _03931_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__xnor2_1
X_06895_ net1069 net1067 net1065 net1072 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__and4bb_4
XANTENNA__08688__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07896__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _03921_ _03922_ _03923_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ cpu.RF0.registers\[1\]\[5\] net713 net709 cpu.RF0.registers\[20\]\[5\] _03845_
+ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout442_A _03594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07516_ net1057 cpu.RF0.registers\[28\]\[6\] net767 vssd1 vssd1 vccd1 vccd1 _02807_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_18_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08496_ cpu.RF0.registers\[6\]\[7\] net675 net635 cpu.RF0.registers\[16\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07112__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08175__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14231__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ net1056 cpu.RF0.registers\[27\]\[1\] net778 vssd1 vssd1 vccd1 vccd1 _02738_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12693__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09839__Y _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08860__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_A _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ cpu.RF0.registers\[20\]\[2\] net594 _02650_ _02654_ _02668_ vssd1 vssd1 vccd1
+ vccd1 _02669_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ _04359_ net291 _04404_ _04394_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a211o_1
XANTENNA__11135__A_N cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14381__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09855__X _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ net1025 cpu.RF0.registers\[20\]\[31\] net780 vssd1 vssd1 vccd1 vccd1 _04339_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07519__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 cpu.RF0.registers\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold471 cpu.RF0.registers\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ cpu.f0.write_data\[25\] _05892_ net993 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__mux2_1
Xhold482 cpu.RF0.registers\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__A2 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 cpu.RF0.registers\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06720__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__A1 cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_1
Xfanout951 _01784_ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_2
Xfanout962 net963 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_2
Xfanout973 net984 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_2
Xfanout984 _01782_ vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_4
XANTENNA__09590__X _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ clknet_leaf_44_clk _00150_ net1305 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13326__Q cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 cpu.RF0.registers\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11772__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1171 cpu.FetchedInstr\[20\] vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 cpu.LCD0.row_2\[31\] vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net2095 net175 net324 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XANTENNA__07887__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ clknet_leaf_29_clk _00023_ net1201 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1193 cpu.RF0.registers\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671__1393 vssd1 vssd1 vccd1 vccd1 _14671__1393/HI net1393 sky130_fd_sc_hd__conb_1
XANTENNA__13329__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__A2 _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14631_ clknet_leaf_31_clk _01732_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11843_ net1631 net209 net330 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14562_ clknet_leaf_51_clk net2472 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_11774_ net1803 net217 net338 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__mux2_1
XANTENNA__07103__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13513_ clknet_leaf_105_clk _00626_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ cpu.IM0.address_IM\[3\] net1015 net286 _05693_ vssd1 vssd1 vccd1 vccd1 _05694_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14493_ clknet_leaf_44_clk _01595_ net1304 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[4\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__13479__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13444_ clknet_leaf_99_clk _00557_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10656_ net2932 cpu.LCD0.row_1\[70\] net907 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XANTENNA__08382__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08813__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload16 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__clkinv_8
X_10587_ net996 net510 _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a21oi_1
Xclkload27 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13375_ clknet_leaf_106_clk _00488_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08603__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__B1 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload38 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload38/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09800__A1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload49 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__clkinv_8
X_12326_ _06202_ net1340 _06201_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__and3b_1
XFILLER_0_23_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__A3 _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ cpu.LCD0.row_1\[86\] _05986_ _06027_ cpu.LCD0.row_2\[46\] _06151_ vssd1 vssd1
+ vccd1 vccd1 _06152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12163__A2 _01965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net1925 net232 net408 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
X_12188_ cpu.LCD0.row_2\[11\] _05998_ _06024_ cpu.LCD0.row_1\[99\] vssd1 vssd1 vccd1
+ vccd1 _06086_ sky130_fd_sc_hd__a22o_1
XANTENNA__10174__A1 cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__B2 cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14620__Q cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ net2781 net249 net416 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
XANTENNA__14104__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06680_ net2270 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[16\] sky130_fd_sc_hd__and2_1
XANTENNA__08557__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14254__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ net943 cpu.RF0.registers\[10\]\[11\] net861 vssd1 vssd1 vccd1 vccd1 _03641_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07301_ cpu.RF0.registers\[1\]\[4\] net589 net571 cpu.RF0.registers\[12\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
X_08281_ net937 cpu.RF0.registers\[11\]\[13\] net880 vssd1 vssd1 vccd1 vccd1 _03572_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07232_ net956 cpu.RF0.registers\[12\]\[9\] net765 vssd1 vssd1 vccd1 vccd1 _02523_
+ sky130_fd_sc_hd__and3_1
XANTENNA_wire877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08723__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07163_ net1043 cpu.RF0.registers\[18\]\[11\] net770 vssd1 vssd1 vccd1 vccd1 _02454_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12018__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07094_ cpu.CU0.funct3\[2\] _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a21o_1
XANTENNA__07339__C net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12139__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11857__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12996__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12154__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07636__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 _05786_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout236 _05770_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
XANTENNA__06908__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09804_ _04496_ _05008_ _05094_ _04480_ _05093_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a221o_1
Xfanout247 _05776_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout269 net271 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ _03284_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or3_1
X_09735_ net299 _04973_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__nand2_1
XANTENNA__12688__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ cpu.RF0.registers\[4\]\[26\] net586 _02216_ _02222_ _02236_ vssd1 vssd1 vccd1
+ vccd1 _02238_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07074__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07869__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _02436_ net300 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__or2_1
X_06878_ net969 net806 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08617_ net1101 cpu.RF0.registers\[30\]\[3\] net840 vssd1 vssd1 vccd1 vccd1 _03908_
+ sky130_fd_sc_hd__and3_1
X_09597_ net301 _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07802__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13621__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08548_ net1107 cpu.RF0.registers\[29\]\[5\] net850 vssd1 vssd1 vccd1 vccd1 _03839_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_59_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ _03766_ _03768_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__or2_1
X_10510_ net1527 net916 net751 a1.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 _00183_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ net1672 net163 net374 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10441_ a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13160_ clknet_leaf_49_clk _00340_ net1376 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[124\]
+ sky130_fd_sc_hd__dfstp_1
X_10372_ a1.curr_state\[0\] net915 _01863_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ net745 _05989_ net557 vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__and3_4
XANTENNA__11767__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ clknet_leaf_53_clk _00271_ net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12452__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14127__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12145__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net556 _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__and2_1
Xhold290 cpu.RF0.registers\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14440__Q cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13151__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout770 _02172_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
Xfanout781 net785 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
Xfanout792 _02150_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
XANTENNA__12598__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ clknet_leaf_2_clk _01106_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07309__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09313__A3 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ clknet_leaf_20_clk _00133_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10459__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06596__S _01965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12875_ clknet_leaf_0_clk cpu.c0.next_count\[6\] net1136 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07712__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11007__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14614_ clknet_leaf_48_clk _01716_ net1362 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[125\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12605__A0 cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ net1900 net147 net336 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__mux2_1
XANTENNA__12869__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ clknet_leaf_50_clk net2187 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_11757_ net2566 net161 net345 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__mux2_1
XANTENNA__08824__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ cpu.LCD0.row_1\[114\] net1680 net897 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ clknet_leaf_33_clk _01586_ net1250 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ net1747 net163 net350 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ clknet_leaf_67_clk _00540_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10639_ cpu.LCD0.row_1\[45\] cpu.LCD0.row_1\[53\] net900 vssd1 vssd1 vccd1 vccd1
+ _00269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_17_clk _00471_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07159__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11677__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ net2866 _01996_ net37 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a21o_1
XANTENNA__10581__S net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12362__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13289_ clknet_leaf_17_clk cpu.RU0.next_FetchedInstr\[28\] net1194 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06998__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10147__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _03137_ _03138_ _03139_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__or4_1
XANTENNA__07563__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _02083_ _02090_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ cpu.RF0.registers\[18\]\[21\] net580 _03050_ _03054_ _03057_ vssd1 vssd1
+ vccd1 vccd1 _03072_ sky130_fd_sc_hd__a2111o_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ _04808_ _04810_ _04801_ _04806_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__o211a_1
XANTENNA__13644__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06732_ net939 net867 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08287__A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07191__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _04739_ _04741_ net486 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__mux2_1
XANTENNA__08718__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06663_ a1.CPU_DAT_O\[31\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07622__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08402_ cpu.RF0.registers\[24\]\[10\] net685 net651 cpu.RF0.registers\[7\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a22o_1
X_09382_ _02348_ _04123_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or2_1
X_06594_ cpu.LCD0.nextState\[3\] net556 _01967_ net1366 vssd1 vssd1 vccd1 vccd1 _01756_
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13794__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ cpu.RF0.registers\[24\]\[12\] net684 net682 cpu.RF0.registers\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09473__C1 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout140_A _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _03545_ _03547_ _03551_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__nor4_1
XFILLER_0_7_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07215_ _02502_ _02504_ _02505_ _02475_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__o31a_1
XANTENNA__13024__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08195_ net1088 cpu.RF0.registers\[26\]\[21\] net860 vssd1 vssd1 vccd1 vccd1 _03486_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10057__A cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ _02436_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08750__A _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07069__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11587__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14670__1392 vssd1 vssd1 vccd1 vccd1 _14670__1392/HI net1392 sky130_fd_sc_hd__conb_1
X_07077_ net1052 cpu.RF0.registers\[29\]\[18\] net793 vssd1 vssd1 vccd1 vccd1 _02368_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13174__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1011 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ net448 _03269_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09718_ net471 _04400_ _04481_ _05007_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__o31a_1
XANTENNA__12296__D1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ cpu.f0.write_data\[19\] _05878_ net990 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07306__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06567__A_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ _03118_ _03402_ _04558_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_2_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12660_ net2126 cpu.LCD0.row_2\[54\] net1005 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__mux2_1
XANTENNA__09059__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ net2241 net201 net359 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08267__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ cpu.IM0.address_IM\[0\] _06350_ _06349_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__mux2_1
X_14330_ clknet_leaf_56_clk _01443_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ net2028 net221 net368 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14261_ clknet_leaf_73_clk _01374_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11473_ net2747 net232 net377 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XANTENNA__09216__C1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07828__X _03119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ clknet_leaf_106_clk _00392_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10424_ net1124 _01817_ net265 vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__or3_1
X_14192_ clknet_leaf_75_clk _01305_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13517__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_53_clk net2624 net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ cpu.f0.i\[27\] _05585_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__or2_1
XANTENNA__08990__A1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ net307 _05525_ _05527_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a31o_1
X_13074_ clknet_leaf_52_clk net2655 net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07707__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12025_ net2192 net142 net313 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__mux2_1
XANTENNA__13667__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10434__C_N cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10430__A cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_6_clk _01089_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12927_ clknet_leaf_26_clk _00116_ net1185 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07442__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11960__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10852__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ clknet_leaf_23_clk _00077_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08835__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08258__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ net1930 net202 net335 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__mux2_1
XANTENNA__13047__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12789_ cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06808__A1 _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528_ clknet_leaf_49_clk _01630_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14459_ clknet_leaf_22_clk _01569_ net1179 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ net1034 cpu.RF0.registers\[16\]\[23\] net831 vssd1 vssd1 vccd1 vccd1 _02291_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13197__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10368__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14442__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08430__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11200__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07186__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ cpu.RF0.registers\[0\]\[27\] net662 net548 vssd1 vssd1 vccd1 vccd1 _04242_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07617__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ cpu.IG0.Instr\[29\] net634 net519 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21o_1
X_08882_ net1080 cpu.RF0.registers\[19\]\[17\] net835 vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14592__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__A2 _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A1 cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ cpu.RF0.registers\[3\]\[24\] net609 net579 cpu.RF0.registers\[18\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a22o_1
XANTENNA__10540__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08729__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10340__A cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ net967 cpu.RF0.registers\[14\]\[21\] net762 vssd1 vssd1 vccd1 vccd1 _03055_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ _03633_ _04051_ net511 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21o_1
X_06715_ net1114 net1110 net1112 net1116 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ net1028 cpu.RF0.registers\[17\]\[17\] net804 vssd1 vssd1 vccd1 vccd1 _02986_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11870__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A _05932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _03019_ net439 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand2_1
X_06646_ a1.CPU_DAT_O\[14\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08745__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09365_ _04522_ _04650_ _02681_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__mux2_1
X_06577_ cpu.K0.count\[0\] cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__nand2_1
XANTENNA_fanout522_A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ net1089 cpu.RF0.registers\[19\]\[12\] net835 vssd1 vssd1 vccd1 vccd1 _03607_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _02213_ _04244_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09461__A2 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_52 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _03534_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10359__A1 cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _03447_ _03452_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__nor3_2
XANTENNA_fanout891_A _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ cpu.RF0.registers\[22\]\[15\] net604 net602 cpu.RF0.registers\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _05405_ _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net626 _04683_ net1023 vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__o21a_1
XANTENNA__10802__X _05749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07527__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_6_clk _00943_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10250__A cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13567__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__A1 cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07262__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ clknet_leaf_63_clk _00874_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10973_ net274 _05865_ _05866_ net926 net2193 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a32o_1
XANTENNA__11780__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10295__B1 cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ net2344 cpu.LCD0.row_2\[106\] net1001 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14315__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13692_ clknet_leaf_8_clk _00805_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12643_ cpu.LCD0.row_2\[45\] cpu.LCD0.row_2\[37\] net997 vssd1 vssd1 vccd1 vccd1
+ _01636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10047__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12574_ cpu.DM0.data_i\[3\] cpu.DM0.data_i\[2\] cpu.DM0.data_i\[5\] cpu.DM0.data_i\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__or4_1
XANTENNA__14465__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14313_ clknet_leaf_104_clk _01426_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ net2546 net179 net371 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__mux2_1
XANTENNA__07463__A1 cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07463__B2 _02753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12907__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14244_ clknet_leaf_98_clk _01357_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11456_ net2160 net167 net381 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
XANTENNA__08390__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06903__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10407_ _01807_ net269 _05621_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11011__A2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14175_ clknet_leaf_0_clk _01288_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ net1762 net188 net387 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13126_ clknet_leaf_54_clk net2565 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ _01893_ _05571_ _05572_ _05574_ net724 vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o311a_1
XANTENNA__07437__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ clknet_leaf_45_clk _00237_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[21\]
+ sky130_fd_sc_hd__dfstp_1
X_10269_ cpu.f0.i\[14\] _05512_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1340 net1341 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_2
X_12008_ net1779 net210 net310 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__mux2_1
Xfanout1351 net1352 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__clkbuf_4
Xfanout1362 net1363 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__clkbuf_2
Xfanout1373 net1377 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__clkbuf_4
Xfanout1384 net1385 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13959_ clknet_leaf_81_clk _01072_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11690__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ _01867_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07480_ net981 cpu.RF0.registers\[13\]\[5\] net794 vssd1 vssd1 vccd1 vccd1 _02771_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09691__A2 _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06431_ cpu.c0.count\[11\] cpu.c0.count\[10\] _01837_ vssd1 vssd1 vccd1 vccd1 _01841_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06362_ cpu.DM0.state\[0\] vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ _04434_ _04440_ net475 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__mux2_1
XANTENNA__10589__A1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ cpu.RF0.registers\[21\]\[22\] net646 net638 cpu.RF0.registers\[26\]\[22\]
+ _03387_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09081_ net460 net447 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _03320_ _03321_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or3_1
XANTENNA__07909__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload42_A clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__C _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold801 cpu.RF0.registers\[28\]\[0\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 cpu.RF0.registers\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 cpu.RF0.registers\[27\]\[13\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 cpu.RF0.registers\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10335__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12026__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 cpu.LCD0.row_2\[79\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 cpu.LCD0.row_2\[115\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 cpu.RF0.registers\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 cpu.RF0.registers\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 cpu.LCD0.row_1\[11\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ net716 net133 _05263_ net629 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a31o_1
XANTENNA__10054__B _05328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ net1084 cpu.RF0.registers\[26\]\[27\] net860 vssd1 vssd1 vccd1 vccd1 _04225_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1501 cpu.LCD0.row_1\[65\] vssd1 vssd1 vccd1 vccd1 net2907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 a1.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1 net2918 sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ _04145_ _04150_ _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout472_A _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1523 cpu.RF0.registers\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net2929 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13212__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14338__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ cpu.RF0.registers\[18\]\[22\] net580 _03084_ _03087_ _03101_ vssd1 vssd1
+ vccd1 vccd1 _03107_ sky130_fd_sc_hd__a2111o_1
X_08796_ _02945_ _03020_ net489 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07390__B1 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12696__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ cpu.RF0.registers\[6\]\[20\] _02175_ _03037_ net623 vssd1 vssd1 vccd1 vccd1
+ _03038_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_101_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07678_ net1024 cpu.RF0.registers\[29\]\[16\] net790 vssd1 vssd1 vccd1 vccd1 _02969_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ _04706_ _04707_ net473 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06629_ _01971_ _01993_ _01994_ _01970_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1267_X net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ _04578_ _04618_ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10229__B cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09279_ net446 net445 net466 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__mux2_1
X_11310_ net2839 net227 net396 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12290_ cpu.LCD0.row_2\[71\] _05988_ _06033_ cpu.LCD0.row_2\[79\] vssd1 vssd1 vccd1
+ vccd1 _06184_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ net1963 net235 net405 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07748__A2 _02160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11172_ net2388 net250 net412 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__mux2_1
XANTENNA__10752__A1 cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13329__Q cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07257__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ cpu.IM0.address_IM\[24\] _03143_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09245__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _05326_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__or2_1
XANTENNA__09370__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08088__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_68_clk _00926_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13705__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ clknet_leaf_75_clk _00857_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10956_ _02543_ net515 _05852_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07133__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13675_ clknet_leaf_89_clk _00788_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ net1804 net207 net430 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13855__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12626_ cpu.LCD0.row_2\[28\] cpu.LCD0.row_2\[20\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12557_ _06309_ _06313_ _01873_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10854__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__X _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__A _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net2778 net224 net371 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__mux2_1
XANTENNA__06633__A a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ net263 _06274_ _06275_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__and3_1
Xhold108 _00155_ vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10991__A1 a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08551__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14623__Q cpu.f0.write_data\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold119 cpu.RF0.registers\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_68_clk _01340_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11439_ net2844 net242 net379 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10155__A cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12193__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07739__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ clknet_leaf_2_clk _01271_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11685__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13235__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ clknet_leaf_51_clk _00289_ net1379 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10442__X _05640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__B _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _02256_ _02258_ _02270_ net619 cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1
+ vccd1 _02271_ sky130_fd_sc_hd__o32ai_4
X_14089_ clknet_leaf_103_clk _01202_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07464__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1170 net1175 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_2
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_4
X_08650_ net1104 cpu.RF0.registers\[18\]\[2\] net853 vssd1 vssd1 vccd1 vccd1 _03941_
+ sky130_fd_sc_hd__and3_1
Xfanout1192 net1199 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13385__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ cpu.RF0.registers\[28\]\[12\] net578 _02873_ _02880_ _02888_ vssd1 vssd1
+ vccd1 vccd1 _02892_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07751__X _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ net1101 cpu.RF0.registers\[25\]\[4\] net863 vssd1 vssd1 vccd1 vccd1 _03872_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14630__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09113__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__B2 _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07470__Y _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ cpu.RF0.registers\[30\]\[6\] _02195_ _02799_ _02805_ _02814_ vssd1 vssd1
+ vccd1 vccd1 _02823_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07463_ cpu.RF0.registers\[0\]\[1\] net618 _02748_ _02753_ vssd1 vssd1 vccd1 vccd1
+ _02754_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_46_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07630__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09202_ _03233_ net434 _04491_ net293 net288 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o221a_1
X_06414_ cpu.c0.count\[6\] cpu.c0.count\[7\] _01826_ vssd1 vssd1 vccd1 vccd1 _01827_
+ sky130_fd_sc_hd__nand3_1
XANTENNA__14277__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07394_ net971 cpu.RF0.registers\[2\]\[0\] net771 vssd1 vssd1 vccd1 vccd1 _02685_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10049__B _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07427__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09133_ net466 _03698_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08624__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout318_A _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09064_ cpu.RF0.registers\[18\]\[31\] net580 _04326_ _04332_ _04346_ vssd1 vssd1
+ vccd1 vccd1 _04355_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_92_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14010__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08461__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ net1097 cpu.RF0.registers\[24\]\[24\] net872 vssd1 vssd1 vccd1 vccd1 _03306_
+ sky130_fd_sc_hd__and3_1
Xhold620 cpu.RF0.registers\[22\]\[15\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 cpu.RF0.registers\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 cpu.RF0.registers\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 cpu.RF0.registers\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07077__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 cpu.RF0.registers\[17\]\[13\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10734__A1 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold675 cpu.RF0.registers\[16\]\[15\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold686 cpu.RF0.registers\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11595__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout687_A _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 cpu.RF0.registers\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _02472_ cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__and2b_1
XANTENNA__14160__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07374__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _04163_ _04198_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__or2_1
XANTENNA__13728__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ cpu.IG0.Instr\[25\] cpu.IM0.address_IM\[5\] net520 vssd1 vssd1 vccd1 vccd1
+ _05185_ sky130_fd_sc_hd__and3_1
XANTENNA__07805__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1320 cpu.LCD0.row_1\[38\] vssd1 vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout854_A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1331 cpu.LCD0.row_1\[73\] vssd1 vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08155__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ net1074 cpu.RF0.registers\[25\]\[16\] net862 vssd1 vssd1 vccd1 vccd1 _04139_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1342 cpu.RF0.registers\[15\]\[12\] vssd1 vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 cpu.LCD0.row_1\[112\] vssd1 vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1364 cpu.RF0.registers\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 cpu.RF0.registers\[4\]\[2\] vssd1 vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 cpu.RF0.registers\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1397 cpu.f0.num\[23\] vssd1 vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ net1100 cpu.RF0.registers\[28\]\[18\] net869 vssd1 vssd1 vccd1 vccd1 _04070_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ net1651 net558 net539 _05754_ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__a22o_1
XANTENNA__13878__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ net1608 net159 net339 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__mux2_1
XANTENNA__07115__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ cpu.f0.data_adr\[8\] _04863_ net993 vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ clknet_leaf_69_clk _00573_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13108__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ net2582 cpu.LCD0.row_1\[86\] net907 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08933__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12411_ cpu.DM0.data_i\[14\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a21o_1
X_13391_ clknet_leaf_86_clk _00504_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12455__A cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07969__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09100__Y _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12342_ _06212_ net1368 _06211_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__and3b_1
XANTENNA__07549__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10973__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14443__Q cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13258__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ _06161_ _06163_ _06165_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__or4_1
XANTENNA__12175__B1 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08918__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14012_ clknet_leaf_12_clk _01125_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ net1892 net167 net407 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
XANTENNA__06740__X _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A1 cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ net1994 net188 net415 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
XANTENNA__13582__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06900__B net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ cpu.IM0.address_IM\[21\] _05355_ cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1
+ vccd1 _05377_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_88_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ cpu.RF0.registers\[2\]\[16\] net205 net422 vssd1 vssd1 vccd1 vccd1 _00520_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07715__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14653__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10037_ cpu.IM0.address_IM\[17\] _02984_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09894__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11988_ net2468 net162 net315 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13727_ clknet_leaf_106_clk _00840_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ net2190 net926 _05675_ net275 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a22o_1
XANTENNA__07450__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13658_ clknet_leaf_86_clk _00771_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14033__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12609_ net2938 cpu.LCD0.row_2\[3\] net997 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XANTENNA__09803__C1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ clknet_leaf_73_clk _00702_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06363__A cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10964__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08281__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14183__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12166__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09031__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09820_ net296 net293 _04930_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__mux2_1
Xfanout407 _05918_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_4
XANTENNA__07465__Y _02756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout418 _05914_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_6
XANTENNA__09393__B _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 _05911_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_4
XANTENNA__07194__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ net479 _04399_ _04631_ _04807_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__o311a_1
X_06963_ cpu.RF0.registers\[22\]\[25\] net604 net569 cpu.RF0.registers\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
XANTENNA__07625__C net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_78_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_08702_ net492 net467 net450 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__or3_1
XANTENNA__08137__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ net487 _03931_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__nand2_1
X_06894_ net962 cpu.RF0.registers\[14\]\[27\] net762 vssd1 vssd1 vccd1 vccd1 _02185_
+ sky130_fd_sc_hd__and3_1
X_08633_ cpu.RF0.registers\[16\]\[3\] net635 _03904_ _03909_ _03910_ vssd1 vssd1 vccd1
+ vccd1 _03924_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12099__X _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout268_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08564_ cpu.RF0.registers\[2\]\[5\] net656 _03839_ _03847_ _03848_ vssd1 vssd1 vccd1
+ vccd1 _03855_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07515_ net978 cpu.RF0.registers\[4\]\[6\] net782 vssd1 vssd1 vccd1 vccd1 _02806_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07360__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08495_ cpu.RF0.registers\[13\]\[7\] net658 net643 cpu.RF0.registers\[3\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ net979 cpu.RF0.registers\[15\]\[1\] net828 vssd1 vssd1 vccd1 vccd1 _02737_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14040__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07377_ net977 cpu.RF0.registers\[14\]\[2\] net763 vssd1 vssd1 vccd1 vccd1 _02668_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13400__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1344_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ _04391_ _04405_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10955__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ net952 cpu.RF0.registers\[14\]\[31\] net761 vssd1 vssd1 vccd1 vccd1 _04338_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12157__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 cpu.RF0.registers\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 cpu.RF0.registers\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10168__C1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 cpu.RF0.registers\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold483 cpu.f0.num\[1\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 cpu.RF0.registers\[24\]\[28\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06720__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_2
X_09949_ cpu.IM0.address_IM\[9\] net933 _05231_ _05232_ vssd1 vssd1 vccd1 vccd1 _00032_
+ sky130_fd_sc_hd__a22o_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_2
Xfanout963 net965 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_69_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net983 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
Xfanout985 net996 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
Xfanout996 cpu.RU0.InstrRead vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_4
X_12960_ clknet_leaf_21_clk _00149_ net1171 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08928__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1150 cpu.RF0.registers\[8\]\[27\] vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__X _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1161 cpu.RF0.registers\[5\]\[1\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net2180 net196 net323 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
Xhold1172 cpu.RF0.registers\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ clknet_leaf_29_clk _00022_ net1201 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1183 cpu.RF0.registers\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 cpu.LCD0.row_1\[71\] vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ clknet_leaf_29_clk _01731_ net1201 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10891__A0 cpu.DM0.readdata\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11842_ net2630 net201 net331 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14056__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14438__Q cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clk_X clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14561_ clknet_leaf_50_clk _01663_ net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ net1632 net221 net340 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__mux2_1
XANTENNA__07270__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13342__Q cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13512_ clknet_leaf_99_clk _00625_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08300__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10724_ cpu.f0.data_adr\[3\] _05030_ net994 vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__mux2_1
X_14492_ clknet_leaf_35_clk _01594_ net1252 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ clknet_leaf_78_clk _00556_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13080__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ cpu.LCD0.row_1\[61\] cpu.LCD0.row_1\[69\] net900 vssd1 vssd1 vccd1 vccd1
+ _00285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload17 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_6
X_13374_ clknet_leaf_86_clk _00487_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10586_ net987 cpu.f0.write_data\[5\] vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nor2_4
XANTENNA__08950__X _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload28 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_6
Xclkload39 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload39/X sky130_fd_sc_hd__clkbuf_8
X_12325_ cpu.LCD0.cnt_20ms\[7\] cpu.LCD0.cnt_20ms\[6\] _05950_ vssd1 vssd1 vccd1 vccd1
+ _06202_ sky130_fd_sc_hd__and3_1
XANTENNA__12148__B1 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_37_clk_X clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__A _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ cpu.LCD0.row_2\[62\] _06000_ _06034_ cpu.LCD0.row_2\[30\] vssd1 vssd1 vccd1
+ vccd1 _06151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11207_ net2701 net244 net408 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
X_12187_ cpu.LCD0.row_2\[3\] _06016_ _06031_ cpu.LCD0.row_1\[27\] _06084_ vssd1 vssd1
+ vccd1 vccd1 _06085_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11138_ net2575 net253 net416 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XANTENNA__07445__C net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09941__B cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _05907_ net503 _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_0_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10579__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13423__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07300_ cpu.RF0.registers\[26\]\[4\] net599 net593 cpu.RF0.registers\[21\]\[4\] _02584_
+ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14549__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ net1082 cpu.RF0.registers\[17\]\[13\] net882 vssd1 vssd1 vccd1 vccd1 _03571_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07231_ net1036 cpu.RF0.registers\[16\]\[9\] net831 vssd1 vssd1 vccd1 vccd1 _02522_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11203__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ net1043 cpu.RF0.registers\[20\]\[11\] net781 vssd1 vssd1 vccd1 vccd1 _02453_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13573__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07093_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06605__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07917__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10343__A cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout204 _05796_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout215 _05793_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
X_09803_ net485 net473 net438 _05008_ net305 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__a311o_1
Xfanout237 _05770_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout248 _05776_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07355__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ cpu.RF0.registers\[1\]\[28\] net713 net709 cpu.RF0.registers\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout385_A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _02604_ _05023_ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__o21a_1
XANTENNA__14639__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__B _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ cpu.RF0.registers\[16\]\[26\] net582 _02215_ _02220_ _02230_ vssd1 vssd1
+ vccd1 vccd1 _02237_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11114__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _04953_ _04954_ _04955_ _04950_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a31o_1
X_06877_ net962 cpu.RF0.registers\[15\]\[27\] net827 vssd1 vssd1 vccd1 vccd1 _02168_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout552_A _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1294_A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ net948 cpu.RF0.registers\[2\]\[3\] net853 vssd1 vssd1 vccd1 vccd1 _03907_
+ sky130_fd_sc_hd__and3_1
X_09596_ _04856_ _04886_ net457 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ cpu.RF0.registers\[10\]\[5\] net693 net635 cpu.RF0.registers\[16\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a22o_1
XANTENNA__08818__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_X net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _03766_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__nand2_1
XANTENNA__12090__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08483__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13916__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07429_ net738 net716 _02092_ net626 _01783_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a41o_2
XFILLER_0_18_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11113__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ a1.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09794__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ _05600_ _05602_ net1590 net729 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12733__A cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10805__X _05751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12940__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _05982_ _05995_ _05996_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_4
X_13090_ clknet_leaf_52_clk _00270_ net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06731__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12452__B cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ net1368 _05950_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__and3_2
XANTENNA__13103__RESET_B net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 cpu.RF0.registers\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 cpu.RF0.registers\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07557__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__B cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _02186_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11783__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 net774 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_8
Xfanout782 net783 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
X_13992_ clknet_leaf_98_clk _01105_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08658__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 _02150_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12302__B1 _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__X _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ clknet_leaf_28_clk _00132_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10313__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ clknet_leaf_0_clk cpu.c0.next_count\[5\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06532__B2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613_ clknet_leaf_49_clk _01715_ net1376 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[124\]
+ sky130_fd_sc_hd__dfstp_1
X_11825_ net2536 net148 net334 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__mux2_1
X_14544_ clknet_leaf_51_clk _01646_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ net2656 net177 net343 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__mux2_1
XANTENNA__07088__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__B1 _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13596__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ cpu.LCD0.row_1\[113\] net1624 net906 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
X_14475_ clknet_leaf_34_clk _01585_ net1251 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10428__A cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ net1636 net167 net351 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__09642__A_N net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12369__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13426_ clknet_leaf_60_clk _00539_ net1344 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10638_ cpu.LCD0.row_1\[44\] cpu.LCD0.row_1\[52\] net904 vssd1 vssd1 vccd1 vccd1
+ _00268_ sky130_fd_sc_hd__mux2_1
XANTENNA__10919__A1 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_102_clk _00470_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10569_ net61 net918 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ net2574 _01996_ net36 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a21o_1
XANTENNA__06641__A a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ clknet_leaf_21_clk cpu.RU0.next_FetchedInstr\[27\] net1173 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[27\] sky130_fd_sc_hd__dfrtp_1
X_12239_ cpu.LCD0.row_1\[85\] _05986_ _06011_ cpu.LCD0.row_2\[53\] _06134_ vssd1 vssd1
+ vccd1 vccd1 _06135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10163__A cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10147__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07012__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14221__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13247__Q a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ _02083_ _02090_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07780_ cpu.RF0.registers\[13\]\[21\] net597 _03047_ _03049_ _03060_ vssd1 vssd1
+ vccd1 vccd1 _03071_ sky130_fd_sc_hd__a2111o_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06731_ net946 net863 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _04698_ _04740_ net471 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__mux2_1
XANTENNA__14371__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06662_ a1.CPU_DAT_O\[30\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[30\]
+ sky130_fd_sc_hd__and2_1
X_08401_ _03678_ _03689_ _03690_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12813__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13939__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ _04582_ _04671_ net481 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06593_ cpu.LCD0.currentState\[3\] net555 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08332_ _03619_ _03620_ _03621_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07079__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload72_A clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08263_ cpu.RF0.registers\[12\]\[15\] net697 _03552_ _03553_ vssd1 vssd1 vccd1 vccd1
+ _03554_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout133_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12963__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07214_ _02493_ _02495_ _02496_ _02497_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ net1084 cpu.RF0.registers\[20\]\[21\] net874 vssd1 vssd1 vccd1 vccd1 _03485_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09225__B1 _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11032__B1 cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07145_ net523 _02433_ _02435_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout300_A _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1042_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13319__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ net1063 cpu.RF0.registers\[26\]\[18\] net788 vssd1 vssd1 vccd1 vccd1 _02367_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07539__A0 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__A cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1307_A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07978_ _03195_ _03197_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10801__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__A _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__inv_2
X_06929_ net1026 cpu.RF0.registers\[22\]\[26\] net799 vssd1 vssd1 vccd1 vccd1 _02220_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07813__C net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11108__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _04936_ _04937_ _04938_ _04927_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_2_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__A4 _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _02581_ _03797_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12599__A0 cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11610_ net2599 net214 net361 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
X_12590_ net630 _05005_ _05149_ _06348_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a22o_1
XANTENNA__06726__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08644__C _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10074__A1 cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net2892 net226 net368 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10248__A cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ clknet_leaf_73_clk _01373_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11472_ net2774 net242 net376 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XANTENNA__07490__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13211_ clknet_leaf_85_clk _00391_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11778__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11023__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _01815_ net269 _05629_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__o21ai_1
X_14191_ clknet_leaf_86_clk _01304_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13142_ clknet_leaf_61_clk _00322_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_10354_ cpu.f0.i\[27\] _05582_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07242__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14244__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14451__Q cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09519__A1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ clknet_leaf_45_clk _00253_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[37\]
+ sky130_fd_sc_hd__dfstp_1
X_10285_ net527 _05528_ _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__and3_1
X_12024_ net2092 net144 net312 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__mux2_1
XANTENNA__14394__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08388__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _02167_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_6
XANTENNA__12836__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ clknet_leaf_66_clk _01088_ net1282 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09152__C1 _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ clknet_leaf_25_clk _00115_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10301__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10857__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ clknet_leaf_23_clk _00076_ net1194 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12986__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ net1696 net212 net335 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__mux2_1
XANTENNA__06636__A a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12788_ net1827 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12357__B net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14626__Q cpu.f0.write_data\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08554__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14527_ clknet_leaf_56_clk net2532 net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_11739_ net2007 net225 net344 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09207__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ clknet_leaf_24_clk _01568_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08851__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11688__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11014__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_63_clk _00522_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09666__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14389_ clknet_leaf_18_clk _01500_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06371__A a1.WRITE_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ net665 _04231_ _04236_ _04240_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__or4b_2
XANTENNA__08981__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13611__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07901_ cpu.RF0.registers\[0\]\[29\] net618 _03188_ _03191_ vssd1 vssd1 vccd1 vccd1
+ _03192_ sky130_fd_sc_hd__o22a_4
XFILLER_0_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08881_ net1077 cpu.RF0.registers\[30\]\[17\] net837 vssd1 vssd1 vccd1 vccd1 _04172_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08733__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _02312_ net259 net488 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_87_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07941__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08729__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ net1039 cpu.RF0.registers\[24\]\[21\] net812 vssd1 vssd1 vccd1 vccd1 _03054_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13761__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ _03633_ _04051_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__nor2_1
X_06714_ _02000_ _02003_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12293__A2 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07694_ net1031 cpu.RF0.registers\[23\]\[17\] net816 vssd1 vssd1 vccd1 vccd1 _02985_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ net484 _04656_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06645_ a1.CPU_DAT_O\[13\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[13\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout250_A _05774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__A _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ net478 _04654_ _04595_ _04535_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__o2bb2a_1
X_06576_ cpu.K0.count\[0\] cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08464__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ net1089 cpu.RF0.registers\[30\]\[12\] net837 vssd1 vssd1 vccd1 vccd1 _03606_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10056__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _02213_ _04244_ net288 vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_42 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1257_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _02410_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09857__A _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13141__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11005__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__B _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _03456_ _03459_ _03463_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or4_1
XANTENNA__06552__Y _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ cpu.RF0.registers\[28\]\[15\] net577 net571 cpu.RF0.registers\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22o_1
XANTENNA__07808__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A _02006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08972__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ cpu.RF0.registers\[0\]\[18\] net618 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__or2_1
XANTENNA__13291__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12859__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ net125 _05343_ _05340_ net626 vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ clknet_leaf_2_clk _00873_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ net987 cpu.f0.write_data\[14\] vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__or2_2
XANTENNA__12284__A2 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08936__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ net2474 net2396 net1005 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__mux2_1
X_13691_ clknet_leaf_13_clk _00804_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12458__A cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12642_ cpu.LCD0.row_2\[44\] cpu.LCD0.row_2\[36\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10047__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14446__Q cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09988__A1 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12573_ _06312_ _06334_ _06335_ _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__o211a_2
XFILLER_0_81_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13350__Q cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14312_ clknet_leaf_84_clk _01425_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11524_ cpu.RF0.registers\[15\]\[23\] net152 net370 vssd1 vssd1 vccd1 vccd1 _00943_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07463__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14243_ clknet_leaf_77_clk _01356_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ net2729 net183 net380 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13634__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ net1126 _01808_ net265 vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__or3_1
X_14174_ clknet_leaf_83_clk _01287_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ net2166 net189 net386 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__mux2_1
X_13125_ clknet_leaf_51_clk _00305_ net1379 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10337_ cpu.f0.i\[24\] _05567_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07574__X _02865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ clknet_leaf_48_clk _00236_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_10268_ cpu.f0.i\[14\] _05512_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13784__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ net1852 net203 net311 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__mux2_1
Xfanout1330 net1331 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1341 net1342 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__buf_2
Xfanout1352 net1356 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__clkbuf_4
X_10199_ _05449_ _05452_ _05460_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__o21ai_1
Xfanout1363 net1364 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__clkbuf_2
Xfanout1374 net1376 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__clkbuf_4
Xfanout1385 net1386 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08549__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11971__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13958_ clknet_leaf_5_clk _01071_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12909_ clknet_leaf_25_clk _00098_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13889_ clknet_leaf_63_clk _01002_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06430_ _01777_ _01838_ _01839_ _01834_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[10\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09428__A0 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06366__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13164__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08284__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__A1 cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08100_ _03384_ _03388_ _03389_ _03390_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_44_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09677__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09080_ _04367_ _04370_ net472 vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07454__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08031_ cpu.RF0.registers\[9\]\[24\] net700 net679 cpu.RF0.registers\[4\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold802 cpu.LCD0.row_2\[89\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09827__D _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11211__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07197__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 cpu.RF0.registers\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07206__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold824 cpu.RF0.registers\[10\]\[4\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 cpu.RF0.registers\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07628__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 cpu.RF0.registers\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload35_A clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold857 cpu.LCD0.row_1\[26\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09982_ cpu.IM0.address_IM\[12\] _05254_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__xor2_1
Xhold868 cpu.RF0.registers\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 cpu.LCD0.row_2\[40\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10761__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net938 cpu.RF0.registers\[14\]\[27\] net838 vssd1 vssd1 vccd1 vccd1 _04224_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14065__RESET_B net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08706__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _04151_ _04152_ _04153_ _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__or4_1
Xhold1502 cpu.RF0.registers\[7\]\[13\] vssd1 vssd1 vccd1 vccd1 net2908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10351__A cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1513 cpu.RF0.registers\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net2919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net2930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1005_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ cpu.RF0.registers\[22\]\[22\] net604 _03092_ _03094_ _03095_ vssd1 vssd1
+ vccd1 vccd1 _03106_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08459__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ cpu.IM0.address_IM\[18\] net553 _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11881__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ cpu.RF0.registers\[14\]\[20\] net575 _02195_ cpu.RF0.registers\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a22o_1
XANTENNA__12266__A2 _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13507__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__B2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07677_ net953 cpu.RF0.registers\[1\]\[16\] net804 vssd1 vssd1 vccd1 vccd1 _02968_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_101_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07142__A1 cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09416_ _04459_ _04469_ net451 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06628_ _01756_ _01976_ _01985_ _01757_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a31o_1
XANTENNA__07693__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _04628_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__nand2_1
X_06559_ net988 _01854_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__nand2_1
XANTENNA__09858__Y _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13657__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ _03371_ _04275_ net460 vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08922__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ cpu.RF0.registers\[27\]\[14\] net712 net652 cpu.RF0.registers\[7\]\[14\]
+ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a221o_1
XANTENNA__06723__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11240_ net2495 net241 net404 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11171_ net2567 net256 net413 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06956__A1 cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ cpu.IM0.address_IM\[23\] net930 _05391_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a21o_1
XANTENNA__08158__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__C1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _05289_ _05300_ _05302_ _05315_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__o41a_2
XANTENNA__10261__A cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ clknet_leaf_69_clk _00925_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06738__X _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__X _04405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10955_ net274 _05853_ _05854_ net926 net2327 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
X_13743_ clknet_leaf_87_clk _00856_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14432__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08330__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ clknet_leaf_101_clk _00787_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07684__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10886_ net723 _05308_ _05808_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a22o_2
XFILLER_0_13_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ net2559 cpu.LCD0.row_2\[19\] net997 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14582__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ _01869_ _06312_ _06310_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_14_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ net2569 net228 net371 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__mux2_1
X_12487_ _05506_ net257 vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07729__B _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06633__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__A2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 cpu.FetchedInstr\[31\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ net1934 net245 net380 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
X_14226_ clknet_leaf_70_clk _01339_ net1326 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07448__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08397__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ clknet_leaf_104_clk _01270_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11369_ net2421 net238 net388 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108_ clknet_leaf_50_clk _00288_ net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ clknet_leaf_98_clk _01201_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ clknet_leaf_44_clk _00219_ net1312 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_37_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__A cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1160 net1162 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_2
Xfanout1171 net1175 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08279__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1182 net1185 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1193 net1199 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
X_07600_ cpu.RF0.registers\[5\]\[12\] net603 _02874_ _02876_ _02883_ vssd1 vssd1 vccd1
+ vccd1 _02891_ sky130_fd_sc_hd__a2111o_1
X_08580_ net1101 cpu.RF0.registers\[22\]\[4\] _02038_ vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12248__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10259__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__S _02756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09113__A2 _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ cpu.RF0.registers\[2\]\[6\] net584 _02802_ _02806_ _02807_ vssd1 vssd1 vccd1
+ vccd1 _02822_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07911__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07462_ _02749_ _02750_ _02751_ _02752_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_46_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09201_ net298 _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__nand2_1
X_06413_ cpu.c0.count\[5\] cpu.c0.count\[4\] _01824_ vssd1 vssd1 vccd1 vccd1 _01826_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07393_ net1048 cpu.RF0.registers\[21\]\[0\] net797 vssd1 vssd1 vccd1 vccd1 _02684_
+ sky130_fd_sc_hd__and3_1
X_09132_ net462 _03664_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07427__A2 _02716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09821__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09200__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ cpu.RF0.registers\[28\]\[31\] net578 _04330_ _04337_ _04338_ vssd1 vssd1
+ vccd1 vccd1 _04354_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload101_A clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ net947 cpu.RF0.registers\[5\]\[24\] net865 vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__and3_1
Xhold610 cpu.RF0.registers\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 cpu.RF0.registers\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07358__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 cpu.DM0.readdata\[31\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 cpu.RF0.registers\[10\]\[11\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 cpu.RF0.registers\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14305__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 cpu.RF0.registers\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 cpu.RF0.registers\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07655__A _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 cpu.RF0.registers\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 cpu.RF0.registers\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09965_ cpu.IM0.address_IM\[11\] _02472_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nand2b_1
X_08916_ _04162_ _04199_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__nor2_1
X_09896_ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__inv_2
Xhold1310 cpu.LCD0.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 cpu.LCD0.row_1\[97\] vssd1 vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08189__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__X _03233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__B2 a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1332 cpu.RF0.registers\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13165__Q a1.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14455__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net1074 cpu.RF0.registers\[20\]\[16\] net874 vssd1 vssd1 vccd1 vccd1 _04138_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07899__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1343 cpu.RF0.registers\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1354 cpu.LCD0.row_2\[86\] vssd1 vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08560__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1365 cpu.RF0.registers\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1376 cpu.RF0.registers\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12239__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1387 cpu.RF0.registers\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ net1100 cpu.RF0.registers\[31\]\[18\] net858 vssd1 vssd1 vccd1 vccd1 _04069_
+ sky130_fd_sc_hd__and3_1
Xhold1398 cpu.RF0.registers\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net2804 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08486__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07729_ _02982_ _03019_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06718__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ net1637 net559 net537 _05704_ vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ cpu.LCD0.row_1\[77\] cpu.LCD0.row_1\[85\] net900 vssd1 vssd1 vccd1 vccd1
+ _00301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12410_ net1615 net732 _06228_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_4_clk _00503_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12411__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__C _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09110__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ cpu.LCD0.cnt_20ms\[13\] cpu.LCD0.cnt_20ms\[12\] _06208_ vssd1 vssd1 vccd1
+ vccd1 _06212_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12272_ cpu.LCD0.row_2\[14\] _05998_ _06011_ cpu.LCD0.row_2\[54\] _06166_ vssd1 vssd1
+ vccd1 vccd1 _06167_ sky130_fd_sc_hd__a221o_1
XANTENNA__07268__C net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ clknet_leaf_11_clk _01124_ net1227 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12175__B2 cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ net2362 net183 net409 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11154_ net2183 net190 net414 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
X_10105_ cpu.IM0.address_IM\[22\] cpu.IM0.address_IM\[21\] _05355_ vssd1 vssd1 vccd1
+ vccd1 _05376_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ net1655 net175 net424 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ cpu.IM0.address_IM\[17\] _02984_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13822__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08827__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ net2746 net180 net317 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__mux2_1
XANTENNA__08303__B1 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ clknet_leaf_84_clk _00839_ net1270 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10938_ net929 cpu.RU0.next_write_i vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__and2b_2
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13972__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ net737 _04813_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__nand2_1
X_13657_ clknet_leaf_92_clk _00770_ net1240 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12608_ cpu.LCD0.row_2\[10\] cpu.LCD0.row_2\[2\] net999 vssd1 vssd1 vccd1 vccd1 _01601_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12402__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06644__A a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_72_clk _00701_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12539_ net1128 cpu.f0.state\[3\] cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 _06307_
+ sky130_fd_sc_hd__nor3_2
XFILLER_0_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13202__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14328__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06890__B_N net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07290__B1 _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11696__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14209_ clknet_leaf_66_clk _01322_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09031__A1 cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13352__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout408 _05918_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_6
Xfanout419 _05914_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09393__C _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ net479 _04625_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o21a_1
X_06962_ cpu.RF0.registers\[24\]\[25\] net608 net599 cpu.RF0.registers\[26\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08701_ cpu.IM0.address_IM\[1\] net553 _03990_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_
+ sky130_fd_sc_hd__a22o_2
X_09681_ net451 _04471_ _03992_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a21bo_1
X_06893_ net966 net764 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08542__B1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ cpu.RF0.registers\[8\]\[3\] net707 net700 cpu.RF0.registers\[9\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a22o_1
XANTENNA__07896__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08563_ cpu.RF0.registers\[7\]\[5\] net653 _03841_ _03844_ net668 vssd1 vssd1 vccd1
+ vccd1 _03854_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07514_ net981 cpu.RF0.registers\[7\]\[6\] net818 vssd1 vssd1 vccd1 vccd1 _02805_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_77_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ cpu.RF0.registers\[4\]\[7\] net678 net667 _03773_ _03780_ vssd1 vssd1 vccd1
+ vccd1 _03785_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_18_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07445_ net979 cpu.RF0.registers\[11\]\[1\] net778 vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout330_A _05938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire809 net810 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_2
X_07376_ net1054 cpu.RF0.registers\[19\]\[2\] net823 vssd1 vssd1 vccd1 vccd1 _02667_
+ sky130_fd_sc_hd__and3_1
X_09115_ _04391_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07288__A2_N net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1337_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ net1026 cpu.RF0.registers\[27\]\[31\] net775 vssd1 vssd1 vccd1 vccd1 _04337_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07820__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 cpu.RF0.registers\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 cpu.RF0.registers\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 cpu.RF0.registers\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 cpu.RF0.registers\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 cpu.RF0.registers\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold495 cpu.RF0.registers\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_2
Xfanout931 _01787_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ _02101_ _04846_ cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o21a_1
Xfanout942 net951 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_2
XANTENNA__13845__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_2
Xfanout975 net983 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_1
Xfanout986 net996 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net1000 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
X_09879_ net125 _05166_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a21o_1
Xhold1140 cpu.RF0.registers\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1151 cpu.LCD0.row_1\[103\] vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 cpu.RF0.registers\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net2229 net198 net325 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
Xhold1173 cpu.RF0.registers\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ clknet_leaf_29_clk _00021_ net1201 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07887__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1184 cpu.RF0.registers\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _00295_ vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09105__A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__A1 _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13995__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__C net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ net2838 net214 net332 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ clknet_leaf_46_clk _01662_ net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07639__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ net2204 net224 net341 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10723_ net1833 net560 net538 _05692_ vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13511_ clknet_leaf_81_clk _00624_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14491_ clknet_leaf_45_clk _01593_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13225__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09111__Y _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ cpu.LCD0.row_1\[60\] cpu.LCD0.row_1\[68\] net904 vssd1 vssd1 vccd1 vccd1
+ _00284_ sky130_fd_sc_hd__mux2_1
X_13442_ clknet_leaf_95_clk _00555_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12185__B _06082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__A1 cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14454__Q cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13373_ clknet_leaf_66_clk _00486_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10585_ _05680_ cpu.LCD0.row_1\[4\] net896 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload18 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_58_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload29 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12324_ cpu.LCD0.cnt_20ms\[6\] _05950_ cpu.LCD0.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ _06201_ sky130_fd_sc_hd__a21o_1
XANTENNA__13375__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__X _02042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ _06111_ _06150_ _06132_ net1354 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__o211a_1
XANTENNA__09494__B _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ net2657 net247 net408 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__07024__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ cpu.LCD0.row_1\[11\] _05994_ _06033_ cpu.LCD0.row_2\[75\] vssd1 vssd1 vccd1
+ vccd1 _06084_ sky130_fd_sc_hd__a22o_1
X_11137_ net1990 net239 net415 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ cpu.IG0.Instr\[7\] cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and2b_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ net627 _05140_ net930 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a21o_1
XANTENNA__07878__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08557__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10882__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13709_ clknet_leaf_102_clk _00822_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14150__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07230_ net956 cpu.RF0.registers\[10\]\[9\] net786 vssd1 vssd1 vccd1 vccd1 _02521_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13718__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12387__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07161_ net966 cpu.RF0.registers\[4\]\[11\] net781 vssd1 vssd1 vccd1 vccd1 _02452_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12387__B2 cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09685__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07092_ net523 _02381_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_67_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13868__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07636__C net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10343__B cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout216 net219 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
X_09802_ _04567_ _04712_ _05091_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a211o_1
Xfanout227 _05786_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 _05770_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
Xfanout249 _05774_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
X_07994_ cpu.RF0.registers\[14\]\[28\] net649 _03273_ _03276_ _03279_ vssd1 vssd1
+ vccd1 vccd1 _03285_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_96_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12892__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _04410_ _04672_ _04680_ _04399_ _04695_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a221o_1
X_06945_ net1026 cpu.RF0.registers\[19\]\[26\] net820 vssd1 vssd1 vccd1 vccd1 _02236_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout280_A _01767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09664_ _03664_ _02473_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__nand2b_1
X_06876_ net972 net830 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__and2_4
XANTENNA__07869__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ net1107 cpu.RF0.registers\[22\]\[3\] _02038_ vssd1 vssd1 vccd1 vccd1 _03906_
+ sky130_fd_sc_hd__and3_1
X_09595_ _04458_ _04468_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__or2_1
XANTENNA__07371__C net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__B _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ _02865_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout712_A _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07428_ cpu.IG0.Instr\[8\] net742 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__nand2_2
XANTENNA__13398__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14643__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ net1054 cpu.RF0.registers\[21\]\[2\] net798 vssd1 vssd1 vccd1 vccd1 _02650_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12573__X _06337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10237__C net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10370_ cpu.f0.i\[29\] _05595_ _05596_ _05601_ net728 vssd1 vssd1 vccd1 vccd1 _05602_
+ sky130_fd_sc_hd__a311o_1
XANTENNA__12733__B _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ _04307_ _04308_ _04318_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__or4_1
XANTENNA__06731__B net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ _05952_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__nor2_1
Xhold270 cpu.RF0.registers\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 cpu.RF0.registers\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07546__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 cpu.RF0.registers\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout750 _05642_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09534__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14023__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_2
X_13991_ clknet_leaf_78_clk _01104_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
Xfanout794 _02150_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08506__B1 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06780__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12942_ clknet_leaf_29_clk _00131_ net1201 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14449__Q cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ clknet_leaf_0_clk cpu.c0.next_count\[4\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13353__Q cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14612_ clknet_leaf_46_clk net1579 net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_11824_ net2540 net155 net334 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__mux2_1
XANTENNA__06746__X _02037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14543_ clknet_leaf_56_clk _01645_ net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09482__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ net2042 net154 net342 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11304__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ cpu.LCD0.row_1\[112\] net1582 net909 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
X_14474_ clknet_leaf_35_clk _01584_ net1251 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_11686_ net2019 net183 net352 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XANTENNA__12369__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__B2 cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13425_ clknet_leaf_76_clk _00538_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net2389 net2407 net899 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10568_ net1133 net1745 net913 _05671_ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13356_ clknet_leaf_67_clk _00469_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08840__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12307_ net2835 net1131 net35 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ net1505 net922 net747 a1.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 _00172_
+ sky130_fd_sc_hd__a22o_1
X_13287_ clknet_leaf_21_clk cpu.RU0.next_FetchedInstr\[26\] net1173 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[26\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06641__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12238_ cpu.LCD0.row_1\[13\] _05994_ _06000_ cpu.LCD0.row_2\[61\] vssd1 vssd1 vccd1
+ vccd1 _06134_ sky130_fd_sc_hd__a22o_1
XANTENNA__11974__S net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__X _05698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ cpu.LCD0.row_2\[66\] _05988_ _06018_ cpu.LCD0.row_2\[98\] _06067_ vssd1 vssd1
+ vccd1 vccd1 _06068_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ net1115 net1113 net1111 net1117 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__and4bb_1
XANTENNA__14516__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06369__A cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10855__A1 _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06661_ a1.CPU_DAT_O\[29\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[29\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07191__C net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ cpu.RF0.registers\[11\]\[10\] net688 _03673_ _03674_ _03680_ vssd1 vssd1
+ vccd1 vccd1 _03691_ sky130_fd_sc_hd__a2111o_1
X_09380_ _04571_ _04670_ net472 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__mux2_1
X_06592_ cpu.LCD0.nextState\[4\] net556 _01966_ net1366 vssd1 vssd1 vccd1 vccd1 _01757_
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08584__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13540__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ cpu.RF0.registers\[27\]\[12\] net711 net708 cpu.RF0.registers\[8\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__a22o_1
XANTENNA__09032__X _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__X _05443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ cpu.RF0.registers\[10\]\[15\] net692 net652 cpu.RF0.registers\[7\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload65_A clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07213_ cpu.RF0.registers\[15\]\[10\] net590 _02503_ net623 vssd1 vssd1 vccd1 vccd1
+ _02504_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08193_ net939 cpu.RF0.registers\[9\]\[21\] net862 vssd1 vssd1 vccd1 vccd1 _03484_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09225__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13690__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ net522 _02434_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07787__A1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__B1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ net973 cpu.RF0.registers\[7\]\[18\] net818 vssd1 vssd1 vccd1 vccd1 _02366_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10354__A cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06551__B _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_98_clk_X clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__A1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__B _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout495_A _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08111__X _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ cpu.IM0.address_IM\[29\] net553 _03266_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_21_clk_X clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14196__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _04594_ _04698_ _04799_ net482 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22oi_2
X_06928_ net954 cpu.RF0.registers\[6\]\[26\] net799 vssd1 vssd1 vccd1 vccd1 _02219_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08197__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ net440 _02348_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__nand2b_1
X_06859_ net1069 net1067 net1065 net1072 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__and4b_4
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _02582_ _03797_ net295 _04868_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08925__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08529_ cpu.RF0.registers\[10\]\[6\] net692 net688 cpu.RF0.registers\[11\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11124__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06726__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ net2080 net228 net368 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XANTENNA__10074__A2 _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ net2856 net246 net376 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
X_10422_ net265 net1124 net1018 vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__or3b_1
X_13210_ clknet_leaf_67_clk _00390_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12220__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09767__A2 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ clknet_leaf_4_clk _01303_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10231__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__A1 cpu.f0.write_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__B2 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ clknet_leaf_52_clk net2728 net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_10353_ _05479_ _05584_ _05587_ net724 cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1
+ _00081_ sky130_fd_sc_hd__o32a_1
XFILLER_0_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10782__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ clknet_leaf_48_clk _00252_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[36\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09519__A2 _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ net541 _05526_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nand2_1
XANTENNA__07276__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__A1 cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net2625 net149 net311 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__mux2_1
XANTENNA__11794__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13413__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14539__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _02179_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_8
Xfanout591 _02165_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_8
XANTENNA__12287__B1 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ clknet_leaf_58_clk _01087_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13563__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ clknet_leaf_26_clk _00114_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14183__RESET_B net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ clknet_leaf_23_clk _00075_ net1194 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ net2576 net218 net334 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__mux2_1
XANTENNA__08258__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12787_ net1444 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06636__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14526_ clknet_leaf_45_clk _01628_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[37\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07466__B1 _02755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ net2518 net228 net344 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11969__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14457_ clknet_leaf_22_clk _01567_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09207__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ net1667 net245 net352 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ clknet_leaf_5_clk _00521_ net1145 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14069__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ clknet_leaf_16_clk _01499_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12762__B2 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__B net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13339_ clknet_leaf_14_clk _00452_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08430__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07186__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13093__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ _03177_ _03180_ _03181_ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__or4_2
XANTENNA__09682__B _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08880_ net1076 cpu.RF0.registers\[21\]\[17\] net866 vssd1 vssd1 vccd1 vccd1 _04171_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08579__A _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07483__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ _02946_ _03021_ _03081_ _02122_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__o31a_1
XANTENNA__07914__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__A1 cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10540__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07762_ net1042 cpu.RF0.registers\[29\]\[21\] net792 vssd1 vssd1 vccd1 vccd1 _03053_
+ sky130_fd_sc_hd__and3_1
X_09501_ net494 _04776_ _04777_ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a31o_2
XFILLER_0_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06713_ _02000_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__and2_4
X_07693_ net1112 _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12930__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ net486 _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__nor2_1
X_06644_ a1.CPU_DAT_O\[12\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06575_ cpu.K0.count\[1\] cpu.K0.count\[0\] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__nand2b_1
X_09363_ _04531_ _04533_ net476 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__mux2_1
XANTENNA__09446__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11253__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ net1089 cpu.RF0.registers\[23\]\[12\] net844 vssd1 vssd1 vccd1 vccd1 _03605_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10056__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09294_ _02213_ _04244_ net293 vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__or3_1
XANTENNA_10 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _02832_ _02868_ _02943_ net490 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a31o_1
XANTENNA__11879__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_43 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__B _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_A _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07658__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ cpu.RF0.registers\[17\]\[20\] net694 _03464_ _03465_ _03466_ vssd1 vssd1
+ vccd1 vccd1 _03467_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08957__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ cpu.RF0.registers\[20\]\[15\] net594 _02415_ _02416_ _02417_ vssd1 vssd1
+ vccd1 vccd1 _02418_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10213__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__B2 cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13436__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09873__A cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ net1111 _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a21o_2
XANTENNA__08709__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__X _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__A2 _02271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08489__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__B1 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _02408_ net516 _05852_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__A _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ net2382 cpu.LCD0.row_2\[104\] net1010 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13690_ clknet_leaf_93_clk _00803_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12458__B cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ net2512 cpu.LCD0.row_2\[35\] net999 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__mux2_1
XANTENNA__09437__A1 _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10047__A2 _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__B1_N net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _01869_ _06311_ _06322_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14211__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ clknet_leaf_82_clk _01424_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11523_ net1872 net164 net370 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14242_ clknet_leaf_96_clk _01355_ net1219 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11454_ net1635 net171 net378 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XANTENNA__14462__Q cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08948__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06903__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net1124 _05620_ net265 net2035 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__a2bb2o_1
X_11385_ net2608 net206 net386 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
X_14173_ clknet_leaf_89_clk _01286_ net1280 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ clknet_leaf_50_clk _00304_ net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09783__A _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10336_ cpu.f0.i\[24\] _05567_ net308 vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13929__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13055_ clknet_leaf_47_clk net2296 net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10267_ _05514_ _05511_ net725 net1547 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1320 net1322 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__clkbuf_4
X_12006_ cpu.RF0.registers\[30\]\[10\] net215 net310 vssd1 vssd1 vccd1 vccd1 _01410_
+ sky130_fd_sc_hd__mux2_1
Xfanout1331 net1342 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__clkbuf_2
Xfanout1342 net1386 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__buf_2
X_10198_ _05449_ _05452_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__or3_1
Xfanout1353 net1355 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__clkbuf_4
Xfanout1364 net1385 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_2
Xfanout1375 net1376 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10522__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1386 net39 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__buf_6
XFILLER_0_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13957_ clknet_leaf_2_clk _01070_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10868__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12908_ clknet_leaf_26_clk _00097_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ clknet_leaf_3_clk _01001_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06647__A a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13309__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12839_ clknet_leaf_30_clk _00058_ net1207 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09428__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06360_ cpu.c0.count\[10\] vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__A2 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11699__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09310__X _04601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ clknet_leaf_47_clk _01611_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09677__B _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08651__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13459__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08030_ cpu.RF0.registers\[16\]\[24\] net637 _03305_ _03314_ _03316_ vssd1 vssd1
+ vccd1 vccd1 _03321_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07478__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07909__C net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold803 _01680_ vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 cpu.LCD0.row_2\[70\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08403__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 cpu.RF0.registers\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10746__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold836 cpu.RF0.registers\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 cpu.LCD0.row_1\[67\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold858 _00250_ vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _05259_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__xor2_1
Xhold869 cpu.RF0.registers\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10903__Y _05822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload28_A clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ net1083 cpu.RF0.registers\[21\]\[27\] net866 vssd1 vssd1 vccd1 vccd1 _04223_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08863_ cpu.RF0.registers\[30\]\[16\] net660 net646 cpu.RF0.registers\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a22o_1
Xhold1503 cpu.RF0.registers\[0\]\[4\] vssd1 vssd1 vccd1 vccd1 net2909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 cpu.f0.num\[4\] vssd1 vssd1 vccd1 vccd1 net2920 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout193_A _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1525 cpu.RF0.registers\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net2931 sky130_fd_sc_hd__dlygate4sd3_1
X_07814_ cpu.RF0.registers\[9\]\[22\] net573 _03097_ _03098_ _03102_ vssd1 vssd1 vccd1
+ vccd1 _03105_ sky130_fd_sc_hd__a2111o_1
X_08794_ cpu.RF0.registers\[0\]\[18\] net663 net549 vssd1 vssd1 vccd1 vccd1 _04085_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12810__RESET_B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07390__A2 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _03029_ _03031_ _03033_ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout360_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07676_ net961 cpu.RF0.registers\[6\]\[16\] net799 vssd1 vssd1 vccd1 vccd1 _02967_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07142__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _04454_ _04461_ net452 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
XANTENNA__14234__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06627_ _01755_ _01985_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06558_ net1130 net1828 net1013 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21o_1
X_09346_ _04415_ _04630_ _04632_ net305 _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__o221a_1
XANTENNA__08772__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09277_ _04427_ _04566_ _04567_ _04441_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06489_ _01876_ _01877_ _01878_ _01879_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__or4_1
XANTENNA__10807__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14384__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08228_ cpu.RF0.registers\[17\]\[14\] net695 net649 cpu.RF0.registers\[14\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout994_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ cpu.RF0.registers\[29\]\[20\] net672 net641 cpu.RF0.registers\[19\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1322_X net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ net2297 net236 net413 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07602__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06956__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net626 _04577_ _05386_ _05390_ net1023 vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o221a_1
XANTENNA__12976__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _05298_ _05313_ _05314_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07554__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__D1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ clknet_leaf_68_clk _00924_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13742_ clknet_leaf_4_clk _00855_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10954_ net986 cpu.f0.write_data\[8\] vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08385__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_104_clk _00786_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ cpu.DM0.readdata\[16\] net734 net719 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__o21a_1
XANTENNA__13601__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ net1584 cpu.LCD0.row_2\[18\] net999 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06754__X _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _01889_ _06309_ _06313_ _01869_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__B1 _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11506_ net2202 net235 net371 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__mux2_1
XANTENNA__07841__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12486_ cpu.f0.i\[11\] net541 net257 cpu.f0.i\[12\] vssd1 vssd1 vccd1 vccd1 _06274_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13751__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ clknet_leaf_77_clk _01338_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ net2865 net251 net380 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10728__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12193__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ clknet_leaf_68_clk _01269_ net1296 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06930__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _05765_ net503 _05920_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__and3_1
XANTENNA__06947__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ clknet_leaf_46_clk net2112 net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _05556_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14107__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ clknet_leaf_80_clk _01200_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11299_ net2812 net143 net401 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ clknet_leaf_45_clk _00218_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11982__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1211 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
Xfanout1172 net1175 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_2
Xfanout1183 net1185 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13131__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__X _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ cpu.RF0.registers\[5\]\[6\] net603 _02804_ _02810_ _02812_ vssd1 vssd1 vccd1
+ vccd1 _02821_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06377__A cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07461_ cpu.RF0.registers\[28\]\[1\] net577 _02727_ _02733_ net623 vssd1 vssd1 vccd1
+ vccd1 _02752_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_46_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13281__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06412_ net1752 _01824_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[4\] sky130_fd_sc_hd__xor2_1
XFILLER_0_31_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09200_ net495 _03234_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07392_ net971 cpu.RF0.registers\[10\]\[0\] net788 vssd1 vssd1 vccd1 vccd1 _02683_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08592__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ _04420_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nor2_1
XANTENNA__08624__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10967__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09062_ cpu.RF0.registers\[5\]\[31\] net603 _04336_ _04340_ _04342_ vssd1 vssd1 vccd1
+ vccd1 _04353_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _03302_ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12999__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold600 cpu.RF0.registers\[29\]\[29\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout206_A _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold611 cpu.RF0.registers\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold622 cpu.RF0.registers\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _01547_ vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 cpu.RF0.registers\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 cpu.RF0.registers\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 cpu.RF0.registers\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06569__B1_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold677 cpu.RF0.registers\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 cpu.RF0.registers\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09964_ cpu.IM0.address_IM\[10\] net933 _05245_ _05246_ vssd1 vssd1 vccd1 vccd1 _00033_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10362__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold699 cpu.RF0.registers\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1115_A cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _03407_ _03442_ _04205_ _03441_ _03405_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__o32a_1
XANTENNA__07374__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ cpu.IG0.Instr\[25\] net520 cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1
+ _05183_ sky130_fd_sc_hd__a21o_1
Xhold1300 _00281_ vssd1 vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11892__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1311 cpu.RF0.registers\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 _00321_ vssd1 vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ net1074 cpu.RF0.registers\[18\]\[16\] net855 vssd1 vssd1 vccd1 vccd1 _04137_
+ sky130_fd_sc_hd__and3_1
Xhold1333 cpu.LCD0.row_1\[96\] vssd1 vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1344 cpu.RF0.registers\[9\]\[25\] vssd1 vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08767__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1355 cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 cpu.RF0.registers\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 cpu.RF0.registers\[8\]\[16\] vssd1 vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ net1100 cpu.RF0.registers\[26\]\[18\] _02025_ vssd1 vssd1 vccd1 vccd1 _04068_
+ sky130_fd_sc_hd__and3_1
Xhold1388 cpu.RF0.registers\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1399 cpu.LCD0.row_1\[72\] vssd1 vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13624__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _02984_ _03018_ net543 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_81_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09731__A1_N _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13181__Q a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ net1024 cpu.RF0.registers\[18\]\[16\] net769 vssd1 vssd1 vccd1 vccd1 _02950_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ cpu.LCD0.row_1\[76\] cpu.LCD0.row_1\[84\] net903 vssd1 vssd1 vccd1 vccd1
+ _00300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08933__C net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13774__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08076__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09329_ _02250_ _04276_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__nor2_1
XANTENNA__10958__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09110__B _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ cpu.LCD0.cnt_20ms\[12\] cpu.LCD0.cnt_20ms\[11\] _06207_ cpu.LCD0.cnt_20ms\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_79_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07549__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10973__A3 _05866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12271_ cpu.LCD0.row_2\[70\] _05988_ _06037_ cpu.LCD0.row_1\[78\] vssd1 vssd1 vccd1
+ vccd1 _06166_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12175__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14010_ clknet_leaf_93_clk _01123_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11222_ net1829 net171 net407 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ net2670 net206 net414 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__mux2_1
XANTENNA__07057__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13154__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net715 net132 _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11084_ net1862 net195 net424 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09879__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ cpu.IM0.address_IM\[16\] net930 _05310_ _05311_ vssd1 vssd1 vccd1 vccd1 _00039_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08000__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11307__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ net2809 net152 net314 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08303__B2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13725_ clknet_leaf_89_clk _00838_ net1280 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10937_ net1802 net131 net430 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__mux2_1
XANTENNA__10110__A1 cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13656_ clknet_leaf_7_clk _00769_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06925__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ net2122 net203 net432 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ net2376 cpu.LCD0.row_2\[1\] net1007 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08067__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13587_ clknet_leaf_68_clk _00700_ net1296 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10799_ net1605 net559 net537 _05746_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a22o_1
XANTENNA__06644__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ net1555 _06304_ _06306_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11977__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10964__A3 _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07290__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ _06262_ _06263_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14208_ clknet_leaf_4_clk _01321_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12166__A2 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06660__A a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10177__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09031__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14139_ clknet_leaf_14_clk _01252_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout409 _05918_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09393__D _04683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09319__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ cpu.RF0.registers\[17\]\[25\] net605 net568 cpu.RF0.registers\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XANTENNA__07194__C net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12323__C1 net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ cpu.RF0.registers\[0\]\[1\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03991_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__13647__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _04969_ _04970_ _04965_ _04967_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12601__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ net1072 net1069 net1067 net1065 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__and4b_1
XANTENNA__07345__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__A1 cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ cpu.RF0.registers\[31\]\[3\] net686 net676 cpu.RF0.registers\[6\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a22o_1
XANTENNA__07922__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ _03838_ _03851_ net542 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13797__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ net1056 cpu.RF0.registers\[17\]\[6\] net806 vssd1 vssd1 vccd1 vccd1 _02804_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ cpu.RF0.registers\[1\]\[7\] net713 _03774_ _03777_ _03778_ vssd1 vssd1 vccd1
+ vccd1 _03784_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10101__A1 cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10101__B2 cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07444_ net1056 cpu.RF0.registers\[20\]\[1\] net782 vssd1 vssd1 vccd1 vccd1 _02735_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ net1054 cpu.RF0.registers\[30\]\[2\] net763 vssd1 vssd1 vccd1 vccd1 _02666_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout323_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _02106_ _02115_ _02116_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__or3b_4
XFILLER_0_33_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09270__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07369__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11887__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A3 _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ net1027 cpu.RF0.registers\[16\]\[31\] net831 vssd1 vssd1 vccd1 vccd1 _04336_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1232_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__A2 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13177__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold430 cpu.RF0.registers\[26\]\[0\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10168__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 cpu.RF0.registers\[19\]\[4\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 a1.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 cpu.RF0.registers\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 cpu.RF0.registers\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 cpu.f0.data_adr\[17\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 cpu.RF0.registers\[25\]\[6\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout910 net911 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_2
Xfanout921 net924 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_5_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09947_ net125 _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_5_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_2
Xfanout954 net961 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net984 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_2
Xfanout976 net978 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_2
Xfanout987 net990 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14572__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ net717 net134 _05167_ net631 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__a31o_1
Xfanout998 net1000 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1130 cpu.RF0.registers\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 cpu.f0.num\[2\] vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 cpu.RF0.registers\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _04114_ _04115_ _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1163 cpu.RF0.registers\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1174 cpu.RF0.registers\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11127__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 cpu.RF0.registers\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 cpu.RF0.registers\[27\]\[7\] vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__B _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11840_ net2578 net218 net330 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08297__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ net2314 net230 net341 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ clknet_leaf_6_clk _00623_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ cpu.IM0.address_IM\[2\] net1015 net285 _05691_ vssd1 vssd1 vccd1 vccd1 _05692_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14490_ clknet_leaf_32_clk _01592_ net1250 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06745__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09121__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ clknet_leaf_63_clk _00554_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ net2431 net2253 net898 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09797__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ clknet_leaf_15_clk _00485_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10584_ net995 _02602_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08960__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload19 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_8
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ _01774_ _05951_ _06200_ net1341 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__o211a_1
XANTENNA__12148__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07576__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ cpu.LCD0.row_1\[125\] _06014_ _06138_ _06140_ _06149_ vssd1 vssd1 vccd1 vccd1
+ _06150_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14137__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06480__A cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ net2855 net251 net409 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XANTENNA__07024__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ net1370 _06082_ _06083_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__and3_1
X_11136_ _05906_ net503 _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__and3_1
XANTENNA__06783__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10730__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net2385 net130 net426 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XANTENNA__09721__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10018_ net125 _05293_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08838__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06639__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11037__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ net2136 net230 net317 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
X_13708_ clknet_leaf_79_clk _00821_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14645__Q cpu.f0.write_data\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ clknet_leaf_82_clk _00752_ net1285 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09788__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07160_ net968 cpu.RF0.registers\[9\]\[11\] net758 vssd1 vssd1 vccd1 vccd1 _02451_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14445__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ net544 _02349_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12139__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07917__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14380__Q cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14595__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 _05810_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_09801_ net272 _04689_ _04708_ _04566_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a22o_1
XANTENNA__07566__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout217 net219 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
XANTENNA__09960__B1 cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
Xfanout239 _05770_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_1
X_07993_ cpu.RF0.registers\[10\]\[28\] net692 net657 cpu.RF0.registers\[13\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkload10_A clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ net481 _04783_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__o21a_1
X_06944_ net1026 cpu.RF0.registers\[26\]\[26\] net786 vssd1 vssd1 vccd1 vccd1 _02235_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09206__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _02508_ _03698_ _04789_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_19_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06875_ net1039 cpu.RF0.registers\[27\]\[27\] net776 vssd1 vssd1 vccd1 vccd1 _02166_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout273_A _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06549__B net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ net1107 cpu.RF0.registers\[25\]\[3\] net863 vssd1 vssd1 vccd1 vccd1 _03905_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06862__A_N net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09594_ _04820_ _04824_ net470 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__mux2_1
X_08545_ _03833_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout440_A _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1182_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10086__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ net491 _02832_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08483__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ net545 _02716_ _02682_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ net976 cpu.RF0.registers\[2\]\[2\] net771 vssd1 vssd1 vccd1 vccd1 _02649_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_18_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07099__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07289_ cpu.IG0.Instr\[27\] net521 net543 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_21_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13812__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ cpu.RF0.registers\[27\]\[31\] net711 net648 cpu.RF0.registers\[25\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 cpu.RF0.registers\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 cpu.RF0.registers\[8\]\[0\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__C1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold282 a1.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07557__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__A2 _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 cpu.RF0.registers\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13962__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 _01853_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_2
Xfanout751 _05642_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
Xfanout762 net764 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_8
X_13990_ clknet_leaf_6_clk _01103_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07309__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__C _02019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08506__B2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ clknet_leaf_29_clk _00130_ net1202 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10313__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__A0 cpu.RF0.registers\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14318__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ clknet_leaf_5_clk cpu.c0.next_count\[3\] net1145 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__A _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ clknet_leaf_54_clk net1535 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[122\]
+ sky130_fd_sc_hd__dfrtp_1
X_11823_ net2011 net159 net335 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14542_ clknet_leaf_45_clk _01644_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[53\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11754_ net2223 net163 net342 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13342__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14468__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10705_ net2402 cpu.LCD0.row_1\[119\] net902 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XANTENNA__14465__Q cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14473_ clknet_leaf_35_clk _01583_ net1250 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08690__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ net1719 net172 net351 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13424_ clknet_leaf_76_clk _00537_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ net2283 net2216 net897 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06762__X _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ clknet_leaf_91_clk _00468_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_10567_ net60 net920 vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__and2_1
XANTENNA__13492__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ net2818 net116 cpu.K0.next_state vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ clknet_leaf_21_clk cpu.RU0.next_FetchedInstr\[25\] net1173 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[25\] sky130_fd_sc_hd__dfrtp_1
X_10498_ net1499 net920 net749 a1.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 _00171_
+ sky130_fd_sc_hd__a22o_1
X_12237_ cpu.LCD0.row_2\[101\] _06018_ _06024_ cpu.LCD0.row_1\[101\] vssd1 vssd1 vccd1
+ vccd1 _06133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ cpu.LCD0.row_1\[90\] _06021_ _06022_ cpu.LCD0.row_2\[122\] vssd1 vssd1 vccd1
+ vccd1 _06067_ sky130_fd_sc_hd__a22o_1
X_11119_ net2863 net205 net418 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
X_12099_ _05982_ _05987_ _05995_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__and3_4
XFILLER_0_78_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07472__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11990__S net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09170__A1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ a1.CPU_DAT_O\[28\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[28\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07720__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06591_ cpu.LCD0.currentState\[4\] _01965_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08330_ cpu.RF0.registers\[11\]\[12\] net690 net656 cpu.RF0.registers\[2\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08261_ cpu.RF0.registers\[6\]\[15\] net675 net635 cpu.RF0.registers\[16\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08681__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13835__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ net1051 cpu.RF0.registers\[31\]\[10\] net830 net566 cpu.RF0.registers\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08192_ net1088 cpu.RF0.registers\[30\]\[21\] net838 vssd1 vssd1 vccd1 vccd1 _03483_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07143_ cpu.IG0.Instr\[15\] _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a21o_1
XANTENNA__08433__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11230__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08984__A1 cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ net974 cpu.RF0.registers\[9\]\[18\] net759 vssd1 vssd1 vccd1 vccd1 _02365_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13985__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1028_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout390_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout488_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13215__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07976_ cpu.RF0.registers\[0\]\[29\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03267_
+ sky130_fd_sc_hd__o21a_1
X_09715_ _04031_ _04033_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__xnor2_1
X_06927_ net958 cpu.RF0.registers\[13\]\[26\] net791 vssd1 vssd1 vccd1 vccd1 _02218_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout655_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _02383_ net441 _04928_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06858_ net963 cpu.RF0.registers\[5\]\[27\] net796 vssd1 vssd1 vccd1 vccd1 _02149_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06847__X _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13365__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _02581_ net436 vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__nor2_1
XANTENNA__14610__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ _02076_ _02077_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout822_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11405__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08528_ cpu.RF0.registers\[1\]\[6\] _02007_ _03804_ _03811_ _03815_ vssd1 vssd1 vccd1
+ vccd1 _03819_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ net1095 cpu.RF0.registers\[25\]\[8\] net863 vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08672__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11470_ net2113 net252 net377 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
X_10421_ net1126 _05628_ net266 net1835 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11023__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08424__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06742__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ clknet_leaf_50_clk _00320_ net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12771__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ _05585_ _05586_ net308 vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_61_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08015__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__A1 a1.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10264__B cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ clknet_leaf_47_clk net2304 net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10283_ cpu.f0.i\[15\] net541 _05518_ cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _05528_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09924__B1 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ net2249 net156 net310 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14140__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _02190_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_8
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08388__C net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout592 _02165_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13708__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ clknet_leaf_69_clk _01086_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12924_ clknet_leaf_25_clk _00113_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12855_ clknet_leaf_39_clk _00074_ net1254 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06917__B _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13858__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ net2032 net220 net336 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ net1421 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14525_ clknet_leaf_48_clk _01627_ net1361 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[36\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07466__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net2357 net234 net344 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__mux2_1
XANTENNA__08663__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09012__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10470__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14456_ clknet_leaf_25_clk _01566_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06492__X _01883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14152__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ net2459 net251 net352 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XANTENNA__06933__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12882__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13407_ clknet_leaf_0_clk _00520_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08851__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ net2516 cpu.LCD0.row_1\[33\] net908 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
XANTENNA__11014__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ clknet_leaf_24_clk _01498_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.CU0.funct3\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11599_ net505 _05907_ _05912_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and3_4
XANTENNA__11050__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12762__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ clknet_leaf_92_clk _00451_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10773__A1 _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11985__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ clknet_leaf_22_clk cpu.RU0.next_FetchedInstr\[8\] net1178 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[8\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09915__B1 cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__X _03503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07830_ _02122_ _03021_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ net1042 cpu.RF0.registers\[26\]\[21\] net787 vssd1 vssd1 vccd1 vccd1 _03052_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14633__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ net278 _04596_ _04779_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a211o_1
X_06712_ cpu.CU0.opcode\[4\] cpu.CU0.opcode\[6\] cpu.CU0.opcode\[3\] cpu.CU0.opcode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__and4b_1
X_07692_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__inv_2
XANTENNA__09694__A2 _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _04720_ _04721_ net475 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06643_ a1.CPU_DAT_O\[11\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[11\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_wire509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11225__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _04482_ _04652_ _04479_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06574_ cpu.K0.count\[0\] cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__or2_1
XANTENNA__09446__A2 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ net1089 cpu.RF0.registers\[28\]\[12\] net869 vssd1 vssd1 vccd1 vccd1 _03604_
+ sky130_fd_sc_hd__and3_1
X_09293_ _02213_ net434 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or2_1
XANTENNA_11 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__X _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout236_A _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__inv_2
XANTENNA_33 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14013__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11005__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ net949 cpu.RF0.registers\[6\]\[20\] net852 vssd1 vssd1 vccd1 vccd1 _03466_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08406__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ net969 cpu.RF0.registers\[8\]\[15\] net813 vssd1 vssd1 vccd1 vccd1 _02417_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07377__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06968__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11895__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__B _02606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07057_ _02315_ _02347_ net543 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_8
XANTENNA_fanout1312_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14163__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__S _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09906__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1100_X net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ net947 cpu.RF0.registers\[10\]\[29\] net861 vssd1 vssd1 vccd1 vccd1 _03250_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12579__X _06342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ net273 _05863_ _05864_ net925 net1952 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a32o_1
XANTENNA__07145__B1 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08936__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _04541_ _04914_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ net2455 cpu.LCD0.row_2\[34\] net999 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09437__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ _06310_ _06313_ _01889_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a21o_1
XANTENNA__12441__A1 cpu.DM0.readdata\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ clknet_leaf_6_clk _01423_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10452__B1 _05640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ net2123 net168 net373 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__mux2_1
XANTENNA__07999__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14241_ clknet_leaf_63_clk _01354_ net1309 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11453_ net2321 net187 net379 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XANTENNA__14506__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ cpu.f0.i\[14\] net269 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__nand2_1
X_14172_ clknet_leaf_11_clk _01285_ net1228 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ net2276 net175 net388 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13123_ clknet_leaf_53_clk _00303_ net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09783__B _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ net1018 cpu.f0.i\[24\] _05560_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07584__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13054_ clknet_leaf_54_clk net2462 net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ net526 _05512_ _05513_ net725 vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13530__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1310 net1313 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09373__A1 _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ net2144 net217 net310 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__mux2_1
Xfanout1321 net1322 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__clkbuf_2
Xfanout1332 net1335 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__clkbuf_4
Xfanout1343 net1364 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__clkbuf_4
X_10197_ _05458_ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1354 net1355 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__clkbuf_4
Xfanout1365 net1367 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__clkbuf_4
Xfanout1376 net1377 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09007__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clk_X clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13680__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07136__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ clknet_leaf_99_clk _01069_ net1232 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06928__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09304__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08846__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ clknet_leaf_25_clk _00096_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13887_ clknet_leaf_0_clk _01000_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11045__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06647__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ clknet_leaf_30_clk _00057_ net1245 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14036__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clk_X clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12769_ net1531 net496 net281 cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14508_ clknet_leaf_46_clk net2832 net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08581__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_clk_X clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13060__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ clknet_leaf_29_clk _01549_ net1188 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10185__A cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14186__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12196__B1 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold804 cpu.RF0.registers\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 cpu.RF0.registers\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07197__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold826 cpu.f0.num\[27\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10746__B2 _05708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 cpu.RF0.registers\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 _00291_ vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12604__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ _05235_ _05238_ _05250_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__o31ai_4
Xhold859 cpu.RF0.registers\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_35_clk_X clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ net1084 cpu.RF0.registers\[28\]\[27\] net869 vssd1 vssd1 vccd1 vccd1 _04222_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12499__B2 cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__B2 _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ cpu.RF0.registers\[1\]\[16\] net714 net670 cpu.RF0.registers\[22\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a22o_1
Xhold1504 cpu.DM0.data_i\[28\] vssd1 vssd1 vccd1 vccd1 net2910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 cpu.RF0.registers\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net2921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 cpu.LCD0.row_1\[62\] vssd1 vssd1 vccd1 vccd1 net2932 sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ net958 cpu.RF0.registers\[6\]\[22\] net800 vssd1 vssd1 vccd1 vccd1 _03104_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12399__X _06223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ _04074_ _04079_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout186_A _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ cpu.RF0.registers\[17\]\[20\] net606 net566 cpu.RF0.registers\[11\]\[20\]
+ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06838__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07660__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ net1024 cpu.RF0.registers\[21\]\[16\] net795 vssd1 vssd1 vccd1 vccd1 _02966_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_101_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout353_A _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ _04697_ _04700_ _04704_ _04694_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a211o_1
X_06626_ _01755_ _01987_ _01992_ _01971_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09501__X _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ net478 _04634_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__o21ai_1
X_06557_ cpu.K0.keyvalid cpu.f0.state\[5\] _01870_ _01942_ vssd1 vssd1 vccd1 vccd1
+ _00023_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout520_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__A cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13403__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14529__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07669__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ net484 _04415_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06488_ cpu.FetchedInstr\[28\] cpu.FetchedInstr\[31\] cpu.FetchedInstr\[30\] cpu.FetchedInstr\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__or4bb_1
XANTENNA__10985__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10985__B2 a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10807__B _04601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ cpu.RF0.registers\[16\]\[14\] net635 _03514_ _03517_ vssd1 vssd1 vccd1 vccd1
+ _03518_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12726__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08158_ cpu.RF0.registers\[15\]\[20\] net683 net657 cpu.RF0.registers\[13\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13179__Q a1.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__X _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ cpu.RF0.registers\[17\]\[14\] net605 net622 vssd1 vssd1 vccd1 vccd1 _02400_
+ sky130_fd_sc_hd__a21o_1
X_08089_ net1086 cpu.RF0.registers\[25\]\[22\] net864 vssd1 vssd1 vccd1 vccd1 _03380_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10120_ net715 net132 _05389_ net627 vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_73_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08158__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12811__Q cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _05324_ _05325_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__nand2_1
XANTENNA__09355__B2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07691__X _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ clknet_leaf_60_clk _00923_ net1344 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12102__X _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ clknet_leaf_104_clk _00854_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10953_ _02864_ net516 _05852_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_67_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08866__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07133__A3 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13672_ clknet_leaf_84_clk _00785_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10884_ net734 net240 vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__nand2_1
XANTENNA__08963__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12623_ net2173 cpu.LCD0.row_2\[17\] net1005 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13083__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07579__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ _06321_ net1641 _06320_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10976__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11505_ net2507 net243 net371 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__mux2_1
X_12485_ _01803_ _06272_ _06273_ net260 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12178__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ clknet_leaf_75_clk _01337_ net1321 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11436_ net2054 net254 net380 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06770__X _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10728__A1 cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08397__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ clknet_leaf_90_clk _01268_ net1278 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11367_ net2535 net129 net390 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__mux2_1
XANTENNA__12920__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_52_clk _00286_ net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10318_ net540 _05556_ _05555_ net526 vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ clknet_leaf_7_clk _01199_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ net2826 net144 net399 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ clknet_leaf_45_clk _00217_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_52_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09346__B2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1151 net1154 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1162 net1167 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10879__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1173 net1175 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1199 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07109__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__A a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14648__Q cpu.f0.write_data\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08857__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13939_ clknet_leaf_67_clk _01052_ net1296 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07480__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_62_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07460_ cpu.RF0.registers\[14\]\[1\] net575 _02721_ _02739_ _02741_ vssd1 vssd1 vccd1
+ vccd1 _02751_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06411_ _01824_ _01825_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[3\] sky130_fd_sc_hd__and2b_1
XFILLER_0_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07391_ cpu.IG0.Instr\[7\] _01851_ _02123_ net1073 vssd1 vssd1 vccd1 vccd1 _02682_
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11503__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ net462 _03729_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14383__Q cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ cpu.RF0.registers\[23\]\[31\] net614 _04331_ _04344_ net621 vssd1 vssd1 vccd1
+ vccd1 _04352_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_96_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ net447 _03301_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload40_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 cpu.RF0.registers\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__B2 cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold612 cpu.RF0.registers\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold623 cpu.RF0.registers\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 cpu.RF0.registers\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 cpu.RF0.registers\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold656 cpu.RF0.registers\[14\]\[26\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 a1.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net632 _04830_ _01787_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 cpu.RF0.registers\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 cpu.RF0.registers\[27\]\[15\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ _03474_ _03510_ _03509_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout1010_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ cpu.IM0.address_IM\[4\] net933 _05181_ _05182_ vssd1 vssd1 vccd1 vccd1 _00027_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10930__X _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1301 cpu.RF0.registers\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ cpu.RF0.registers\[12\]\[16\] net696 _04133_ _04134_ _04135_ vssd1 vssd1
+ vccd1 vccd1 _04136_ sky130_fd_sc_hd__a2111o_1
Xhold1312 cpu.RF0.registers\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 cpu.RF0.registers\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14201__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1334 cpu.RF0.registers\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 cpu.RF0.registers\[21\]\[23\] vssd1 vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout568_A _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1356 cpu.LCD0.row_1\[22\] vssd1 vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 cpu.RF0.registers\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ net948 cpu.RF0.registers\[2\]\[18\] net853 vssd1 vssd1 vccd1 vccd1 _04067_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06571__A1 cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1378 cpu.RF0.registers\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 cpu.RF0.registers\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08486__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07727_ cpu.RF0.registers\[0\]\[17\] net617 _03014_ _03017_ vssd1 vssd1 vccd1 vccd1
+ _03018_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_81_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14351__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ net953 cpu.RF0.registers\[15\]\[16\] net825 vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06855__X _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13919__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06609_ _01974_ _01755_ _01978_ _01971_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout902_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07589_ net1046 cpu.RF0.registers\[19\]\[12\] net821 vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11413__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09328_ _02250_ _04276_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_24_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10537__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12806__Q cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09259_ _04414_ _04537_ _04545_ _04480_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12943__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ cpu.LCD0.row_1\[38\] _06006_ _06031_ cpu.LCD0.row_1\[30\] _06164_ vssd1 vssd1
+ vccd1 vccd1 _06165_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09025__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06590__X _01965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11221_ cpu.RF0.registers\[6\]\[18\] net187 net408 vssd1 vssd1 vccd1 vccd1 _00650_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11152_ net2284 net175 net416 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
XANTENNA__08023__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _05371_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__xnor2_1
X_11083_ net2793 net198 net425 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08958__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10034_ net627 net240 net930 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13449__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11985_ net1795 net163 net314 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09500__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13724_ clknet_leaf_8_clk _00837_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ _05474_ _05844_ net719 vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13599__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ net722 _05256_ _05794_ _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13655_ clknet_leaf_66_clk _00768_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11323__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ net2349 cpu.LCD0.row_2\[0\] net1008 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13586_ clknet_leaf_60_clk _00699_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ cpu.IM0.address_IM\[24\] net1014 net285 _05745_ vssd1 vssd1 vccd1 vccd1 _05746_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__Y _05086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ cpu.f0.i\[31\] _06304_ net260 vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07290__A2 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12468_ cpu.f0.i\[5\] _06260_ net261 vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09016__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06941__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14207_ clknet_leaf_106_clk _01320_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11419_ net2182 net191 net382 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12399_ cpu.DM0.data_i\[8\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07578__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06660__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10177__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14138_ clknet_leaf_94_clk _01251_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14224__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07475__C net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09319__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ net1044 cpu.RF0.registers\[23\]\[25\] net817 vssd1 vssd1 vccd1 vccd1 _02251_
+ sky130_fd_sc_hd__and3_1
X_14069_ clknet_leaf_73_clk _01182_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_3_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11126__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06891_ net1050 net767 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__and2_2
XFILLER_0_94_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08630_ cpu.RF0.registers\[10\]\[3\] net693 _03905_ _03913_ _03914_ vssd1 vssd1 vccd1
+ vccd1 _03921_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08542__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14374__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06553__A1 cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08561_ cpu.RF0.registers\[9\]\[5\] net700 _03843_ _03846_ _03850_ vssd1 vssd1 vccd1
+ vccd1 _03852_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07512_ net981 cpu.RF0.registers\[14\]\[6\] net764 vssd1 vssd1 vccd1 vccd1 _02803_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08492_ cpu.RF0.registers\[7\]\[7\] net652 _03772_ _03781_ _03782_ vssd1 vssd1 vccd1
+ vccd1 _03783_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10101__A2 _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload88_A clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07443_ net979 cpu.RF0.registers\[4\]\[1\] net782 vssd1 vssd1 vccd1 vccd1 _02734_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12966__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ net979 cpu.RF0.registers\[15\]\[2\] net828 vssd1 vssd1 vccd1 vccd1 _02665_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09113_ net437 _04399_ _04402_ _04358_ _04398_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08463__D1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout316_A _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1058_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ net961 cpu.RF0.registers\[8\]\[31\] net811 vssd1 vssd1 vccd1 vccd1 _04335_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07281__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 cpu.DM0.readdata\[21\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 cpu.RF0.registers\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06570__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 cpu.RF0.registers\[1\]\[29\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1225_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 cpu.FetchedInstr\[11\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 cpu.RF0.registers\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 cpu.DM0.readdata\[10\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 cpu.RF0.registers\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout685_A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout911 _01940_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
Xhold497 cpu.RF0.registers\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08781__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ net717 net134 _05229_ net631 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 _01787_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14436__RESET_B net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_2
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_2
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_1
Xhold1120 cpu.LCD0.row_1\[115\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ cpu.IM0.address_IM\[3\] cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 _05167_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout852_A _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net990 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1131 cpu.RF0.registers\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11408__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1142 cpu.RF0.registers\[5\]\[12\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 cpu.LCD0.row_2\[27\] vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ cpu.RF0.registers\[15\]\[19\] net683 _04116_ _04117_ _04118_ vssd1 vssd1
+ vccd1 vccd1 _04119_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_68_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 cpu.RF0.registers\[18\]\[21\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 a1.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 cpu.RF0.registers\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _04043_ _04046_ _04048_ _03669_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1197 cpu.RF0.registers\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13741__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11770_ net1830 net233 net340 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10721_ cpu.f0.data_adr\[2\] _05043_ net992 vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06745__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13891__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ clknet_leaf_3_clk _00553_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10652_ net2433 net1805 net902 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__mux2_1
XANTENNA__09246__A0 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08018__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13371_ clknet_leaf_12_clk _00484_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10583_ net987 cpu.f0.write_data\[4\] vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_58_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ _01774_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__nand2_1
XANTENNA__13121__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14247__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ _06142_ _06144_ _06146_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__or4_1
XANTENNA__07576__B _02865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06480__B _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__A2 _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ net2523 net254 net409 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__mux2_1
XANTENNA__07024__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ net121 net555 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__or2_1
XANTENNA__13271__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ cpu.IG0.Instr\[10\] cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__and2b_2
XFILLER_0_21_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14397__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ net2237 net136 net426 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XANTENNA__10730__B _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net715 net132 _05294_ net627 vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07732__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__A1 cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12989__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06936__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ cpu.RF0.registers\[29\]\[5\] net233 net316 vssd1 vssd1 vccd1 vccd1 _01373_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10095__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ clknet_leaf_91_clk _00820_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ cpu.DM0.readdata\[26\] _04640_ net734 vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11899_ net1838 net249 net323 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
XANTENNA__11053__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13638_ clknet_leaf_5_clk _00751_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09788__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__S net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09966__B cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10892__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__X _05708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13569_ clknet_leaf_66_clk _00682_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ _02377_ _02379_ _02380_ _02350_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__o31a_2
XFILLER_0_67_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10905__B _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13614__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__A cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09960__A1 cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ net291 _05089_ _05090_ net444 _03045_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__o32a_1
Xfanout207 _05810_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
X_07992_ net1093 cpu.RF0.registers\[24\]\[28\] net871 vssd1 vssd1 vccd1 vccd1 _03283_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _04384_ _04875_ _05021_ _02759_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__o2bb2a_1
X_06943_ net1026 cpu.RF0.registers\[25\]\[26\] net756 vssd1 vssd1 vccd1 vccd1 _02234_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13764__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _04789_ _04951_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__or3_1
X_06874_ net1050 net777 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__and2_1
X_08613_ net1107 cpu.RF0.registers\[29\]\[3\] net850 vssd1 vssd1 vccd1 vccd1 _03904_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09593_ _04607_ _04883_ _04807_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ _02830_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06846__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10086__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ _03764_ _03765_ cpu.IM0.address_IM\[8\] net554 vssd1 vssd1 vccd1 vccd1 _03766_
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1175_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ net545 _02716_ _02682_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13144__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07357_ net976 cpu.RF0.registers\[8\]\[2\] net813 vssd1 vssd1 vccd1 vccd1 _02648_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout600_A _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1342_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ cpu.RF0.registers\[0\]\[7\] net618 net518 net517 vssd1 vssd1 vccd1 vccd1
+ _02579_ sky130_fd_sc_hd__a2bb2o_4
X_09027_ cpu.RF0.registers\[23\]\[31\] net671 net670 cpu.RF0.registers\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13294__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1130_X net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1228_X net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 cpu.RF0.registers\[12\]\[10\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 cpu.RF0.registers\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13187__Q a1.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 cpu.RF0.registers\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A1 cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 cpu.RF0.registers\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 cpu.RF0.registers\[29\]\[10\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 net732 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_2
XANTENNA__07962__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout752 _05639_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
X_09929_ cpu.IM0.address_IM\[8\] _02833_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__xnor2_1
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11138__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout796 net798 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
X_12940_ clknet_leaf_29_clk _00129_ net1202 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09116__B _04405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ clknet_leaf_5_clk cpu.c0.next_count\[2\] net1145 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[2\] sky130_fd_sc_hd__dfrtp_1
X_14610_ clknet_leaf_52_clk net1492 net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12110__X _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ net2464 net179 net336 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14541_ clknet_leaf_48_clk _01643_ net1361 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_11753_ net1657 net168 net345 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ net2429 net2493 net908 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
X_14472_ clknet_leaf_35_clk _01582_ net1251 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07493__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11684_ net2611 net188 net352 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11026__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10635_ net2365 cpu.LCD0.row_1\[49\] net906 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
X_13423_ clknet_leaf_81_clk _00536_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12493__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ clknet_leaf_95_clk _00467_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07587__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ net1134 net1651 net914 _05670_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__a31o_1
XANTENNA__07245__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14481__Q a1.WRITE_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ cpu.K0.code\[2\] net115 cpu.K0.next_state vssd1 vssd1 vccd1 vccd1 _01458_
+ sky130_fd_sc_hd__mux2_1
X_13285_ clknet_leaf_21_clk cpu.RU0.next_FetchedInstr\[24\] net1173 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[24\] sky130_fd_sc_hd__dfrtp_1
X_10497_ net82 net922 net747 net1425 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236_ net2928 net555 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10001__A1 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ cpu.LCD0.row_1\[82\] _05986_ _06015_ cpu.LCD0.row_1\[2\] _06065_ vssd1 vssd1
+ vccd1 vccd1 _06066_ sky130_fd_sc_hd__a221o_1
X_11118_ net2010 net173 net420 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__mux2_1
X_12098_ cpu.LCD0.row_1\[8\] _05994_ _05998_ cpu.LCD0.row_2\[8\] vssd1 vssd1 vccd1
+ vccd1 _05999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13017__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11048__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ net2089 net197 net426 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__mux2_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09170__A2 _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10887__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06913__D1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06590_ _01956_ _01962_ _01963_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__and4bb_2
XANTENNA__06666__A a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08584__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__A1 cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14412__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08130__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _03542_ _03548_ _03549_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08881__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07211_ _02498_ _02499_ _02500_ _02501_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__or4_1
XANTENNA__11017__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08191_ net1088 cpu.RF0.registers\[31\]\[21\] net859 vssd1 vssd1 vccd1 vccd1 _03482_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12765__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14562__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ cpu.RF0.registers\[0\]\[15\] net619 _02422_ _02432_ vssd1 vssd1 vccd1 vccd1
+ _02433_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_67_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06832__C net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14391__Q cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ net1052 cpu.RF0.registers\[22\]\[18\] net803 vssd1 vssd1 vccd1 vccd1 _02364_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08984__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09933__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07663__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ net667 _03256_ _03261_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout383_A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ _04911_ _05004_ _04904_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__or3b_4
X_06926_ net1026 cpu.RF0.registers\[24\]\[26\] net811 vssd1 vssd1 vccd1 vccd1 _02217_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12296__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09645_ _04932_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nand2_1
XANTENNA__10797__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06857_ net967 net796 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout550_A _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1292_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ _02582_ _03797_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06788_ cpu.RF0.registers\[12\]\[30\] net696 net636 cpu.RF0.registers\[16\]\[30\]
+ _02046_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a221o_1
XANTENNA__14092__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ cpu.RF0.registers\[27\]\[6\] net712 net647 cpu.RF0.registers\[21\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__A cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ net946 cpu.RF0.registers\[11\]\[8\] net879 vssd1 vssd1 vccd1 vccd1 _03749_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06863__X _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__A1 cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11008__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07409_ net1048 cpu.RF0.registers\[17\]\[0\] net806 vssd1 vssd1 vccd1 vccd1 _02700_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08389_ net945 cpu.RF0.registers\[4\]\[10\] net877 vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10826__A cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net1019 net270 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__nand2_1
XANTENNA__12213__B1_N net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12220__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12814__Q cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07200__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ cpu.f0.i\[26\] _05579_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__nand2_1
XANTENNA__08975__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__B1 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10782__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ clknet_leaf_54_clk net2264 net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__inv_2
X_12021_ net1884 net161 net312 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__A1 cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12105__X _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
Xfanout571 net572 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_8
Xfanout582 _02177_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_8
XANTENNA__12287__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout593 _02162_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_8
X_13972_ clknet_leaf_69_clk _01085_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08966__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A1 cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__X _04705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ clknet_leaf_22_clk _00112_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14435__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12854_ clknet_leaf_38_clk _00073_ net1262 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11805_ net2240 net226 net337 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__mux2_1
X_12785_ net1511 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14585__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ clknet_leaf_46_clk _01626_ net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__A2 _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__X _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11736_ net2618 net244 net344 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14455_ clknet_leaf_25_clk _01565_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10470__B2 a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net1893 net255 net353 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11331__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__B1 _06345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13406_ clknet_leaf_85_clk _00519_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ net2617 net2226 net909 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
X_14386_ clknet_leaf_24_clk _01497_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.CU0.funct3\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11598_ net1739 net128 net362 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XANTENNA__10222__A1 cpu.f0.data_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ net50 net921 vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__and2_1
XANTENNA__10222__B2 cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13337_ clknet_leaf_42_clk _00450_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13268_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[7\] net1246 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[7\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_47_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08179__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A1 _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ cpu.LCD0.row_2\[4\] _06016_ _06019_ cpu.LCD0.row_1\[52\] _06115_ vssd1 vssd1
+ vccd1 vccd1 _06116_ sky130_fd_sc_hd__a221o_1
X_13199_ clknet_leaf_70_clk _00379_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07483__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07760_ net1042 cpu.RF0.registers\[25\]\[21\] net757 vssd1 vssd1 vccd1 vccd1 _03051_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12278__A2 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ _01999_ _02000_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__nand2_2
X_07691_ _02947_ _02981_ net543 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_4
XFILLER_0_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09430_ _04570_ _04668_ net455 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__mux2_1
XANTENNA__11506__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06642_ a1.CPU_DAT_O\[10\] net895 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[10\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__13802__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06396__A cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14386__Q cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ net479 _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nand2_1
X_06573_ _01833_ cpu.c0.next_count\[16\] _01952_ cpu.c0.next_count\[0\] vssd1 vssd1
+ vccd1 vccd1 cpu.c0.next_atmax sky130_fd_sc_hd__and4b_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09446__A3 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08312_ cpu.RF0.registers\[12\]\[12\] net698 net659 cpu.RF0.registers\[13\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a22o_1
XANTENNA__09300__C1 _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ _04412_ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_9_clk_X clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload70_A clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13952__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ cpu.IM0.address_IM\[14\] net553 _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__a22o_4
XANTENNA_34 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ net1099 cpu.RF0.registers\[24\]\[20\] net872 vssd1 vssd1 vccd1 vccd1 _03465_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07209__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ net1050 cpu.RF0.registers\[29\]\[15\] net793 vssd1 vssd1 vccd1 vccd1 _02416_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08957__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10933__X _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14308__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10764__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07955__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _02342_ _02344_ _02346_ _02316_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09906__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1305_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08489__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14458__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__X _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ net1097 cpu.RF0.registers\[23\]\[29\] net845 vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__and3_1
X_06909_ cpu.RF0.registers\[28\]\[27\] net578 _02185_ _02168_ _02176_ vssd1 vssd1
+ vccd1 vccd1 _02200_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07145__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07889_ cpu.RF0.registers\[16\]\[29\] net581 net574 cpu.RF0.registers\[9\]\[29\]
+ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13482__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _03172_ net447 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__xor2_1
XANTENNA__12809__Q cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _04848_ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12570_ _01867_ _06311_ _06313_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ net2659 net183 net371 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10452__B2 a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11151__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ net1840 net189 net378 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
X_14240_ clknet_leaf_2_clk _01353_ net1154 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08026__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ net1125 _05619_ net264 net2129 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10204__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08948__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14171_ clknet_leaf_14_clk _01284_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10990__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ net2353 net193 net388 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__mux2_1
XANTENNA__06959__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ clknet_leaf_56_clk net2583 net1371 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_10334_ net1018 _05560_ cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13053_ clknet_leaf_52_clk net2131 net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10265_ cpu.f0.i\[13\] _05506_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__nor2_1
Xfanout1300 net1386 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__clkbuf_4
X_12004_ net2014 net223 net312 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__mux2_1
Xfanout1311 net1313 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_2
XFILLER_0_24_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1322 net1342 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_2
X_10196_ cpu.IM0.address_IM\[30\] _03232_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__or2_1
Xfanout1333 net1334 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__clkbuf_4
Xfanout1344 net1364 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__clkbuf_2
Xfanout1355 net1356 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__buf_2
Xfanout1366 net1367 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13825__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1377 net1385 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_92_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06768__X _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout390 net393 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13955_ clknet_leaf_77_clk _01068_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11326__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ clknet_leaf_26_clk _00095_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload7_A clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__B net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ clknet_leaf_85_clk _00999_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13975__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12837_ clknet_leaf_30_clk _00056_ net1208 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06944__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12768_ net1539 net496 net281 cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14507_ clknet_leaf_54_clk _01609_ net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11719_ net2348 net181 net347 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12699_ cpu.LCD0.row_2\[101\] cpu.LCD0.row_2\[93\] net998 vssd1 vssd1 vccd1 vccd1
+ _01692_ sky130_fd_sc_hd__mux2_1
XANTENNA__11061__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06663__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14438_ clknet_leaf_29_clk _01548_ net1189 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14302__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__C net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11996__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08939__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14369_ clknet_leaf_27_clk cpu.K0.next_state net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.state
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold805 cpu.f0.num\[25\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 cpu.RF0.registers\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10746__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold827 cpu.LCD0.row_2\[46\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 cpu.RF0.registers\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13355__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 cpu.RF0.registers\[0\]\[29\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14600__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08930_ net1084 cpu.RF0.registers\[25\]\[27\] net862 vssd1 vssd1 vccd1 vccd1 _04221_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ cpu.RF0.registers\[4\]\[16\] net677 net638 cpu.RF0.registers\[26\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__a22o_1
Xhold1505 cpu.RF0.registers\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net2911 sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ net1032 cpu.RF0.registers\[27\]\[22\] net776 vssd1 vssd1 vccd1 vccd1 _03103_
+ sky130_fd_sc_hd__and3_1
Xhold1516 cpu.LCD0.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 a1.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net2933 sky130_fd_sc_hd__dlygate4sd3_1
X_08792_ _04061_ _04080_ _04081_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or4_1
XFILLER_0_93_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07743_ cpu.RF0.registers\[19\]\[20\] net615 net570 cpu.RF0.registers\[10\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08324__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06838__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07674_ net1024 cpu.RF0.registers\[24\]\[16\] net811 vssd1 vssd1 vccd1 vccd1 _02965_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_101_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09783__D_N _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ _04702_ _04703_ _03173_ net447 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__o2bb2a_1
X_06625_ _01972_ _01974_ _01981_ _01970_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout346_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06556_ _01780_ cpu.f0.state\[7\] vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _04385_ _04503_ _04633_ _04382_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o211a_1
XANTENNA__08772__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ net478 _04383_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__A cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06487_ cpu.FetchedInstr\[25\] cpu.FetchedInstr\[24\] cpu.FetchedInstr\[27\] cpu.FetchedInstr\[26\]
+ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1255_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08226_ cpu.RF0.registers\[31\]\[14\] net686 _03515_ _03516_ vssd1 vssd1 vccd1 vccd1
+ _03517_ sky130_fd_sc_hd__a211o_1
XANTENNA__14043__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12187__A1 cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ cpu.RF0.registers\[12\]\[20\] net697 net648 cpu.RF0.registers\[25\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07108_ cpu.RF0.registers\[1\]\[14\] net588 net568 cpu.RF0.registers\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a22o_1
XANTENNA__11034__A_N cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08088_ net1080 cpu.RF0.registers\[22\]\[22\] net851 vssd1 vssd1 vccd1 vccd1 _03379_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07602__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14280__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07039_ net963 cpu.RF0.registers\[6\]\[19\] _02145_ vssd1 vssd1 vccd1 vccd1 _02330_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1210_X net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13848__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10050_ cpu.IM0.address_IM\[18\] _02349_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13998__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06748__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_80_clk _00853_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10952_ net992 _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nand2_4
XANTENNA__08866__A1 cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ clknet_leaf_80_clk _00784_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10883_ net2027 net176 net432 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
X_12622_ net2412 net2194 net1007 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06764__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ net1128 cpu.DM0.data_i\[0\] _06307_ _06316_ vssd1 vssd1 vccd1 vccd1 _06321_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09291__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__A2 cpu.f0.write_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11504_ net1928 net245 net371 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _01803_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__nand2_1
XANTENNA__07841__A2 _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13378__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ clknet_leaf_82_clk _01336_ net1285 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11435_ net2108 net238 net379 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07054__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07595__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14154_ clknet_leaf_102_clk _01267_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11366_ net1567 net138 net390 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__mux2_1
XANTENNA__06930__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13105_ clknet_leaf_48_clk _00285_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[69\]
+ sky130_fd_sc_hd__dfstp_1
X_10317_ cpu.f0.i\[21\] _05549_ net307 vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ net2556 net150 net399 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
X_14085_ clknet_leaf_9_clk _01198_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ clknet_leaf_45_clk _00216_ net1312 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_10248_ cpu.f0.i\[11\] _05491_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1130 a1.BUSY_O vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_2
XFILLER_0_20_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1141 net1143 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1152 net1154 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ cpu.IM0.address_IM\[27\] _05422_ cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1
+ vccd1 _05444_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10361__B1 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1163 net1166 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1174 net1175 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_2
Xfanout1185 net1191 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XANTENNA__14003__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07761__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1196 net1198 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11056__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13938_ clknet_leaf_60_clk _01051_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13869_ clknet_leaf_105_clk _00982_ net1156 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14153__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06410_ cpu.c0.count\[1\] cpu.c0.count\[0\] cpu.c0.count\[2\] cpu.c0.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ net524 _02679_ _02645_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o21ai_4
XANTENNA__06674__A a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12405__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08592__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09060_ _04347_ _04348_ _04349_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_96_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07293__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ net447 _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__and2_1
XANTENNA__07001__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10719__A2 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold602 cpu.RF0.registers\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11916__A1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 cpu.RF0.registers\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 cpu.RF0.registers\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 cpu.RF0.registers\[17\]\[27\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload33_A clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold646 cpu.LCD0.row_1\[31\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 cpu.RF0.registers\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 cpu.f0.num\[0\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 a1.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net127 _05244_ _05241_ net632 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08913_ _04055_ _04056_ _04202_ _03513_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a211o_1
XANTENNA__12895__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ net625 _05016_ net1022 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 cpu.RF0.registers\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ net1074 cpu.RF0.registers\[23\]\[16\] net844 vssd1 vssd1 vccd1 vccd1 _04135_
+ sky130_fd_sc_hd__and3_1
Xhold1313 cpu.RF0.registers\[7\]\[7\] vssd1 vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07899__A2 _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06849__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 cpu.RF0.registers\[1\]\[25\] vssd1 vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 cpu.RF0.registers\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 cpu.DM0.readdata\[2\] vssd1 vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08767__C _02019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1357 cpu.RF0.registers\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07671__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1368 cpu.RF0.registers\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ net1109 cpu.RF0.registers\[21\]\[18\] net865 vssd1 vssd1 vccd1 vccd1 _04066_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1379 cpu.K0.code\[7\] vssd1 vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
X_07726_ _03008_ _03009_ _03015_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_81_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ net953 cpu.RF0.registers\[14\]\[16\] net761 vssd1 vssd1 vccd1 vccd1 _02948_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14295__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06608_ _01974_ _01977_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nand2_1
X_07588_ net1045 cpu.RF0.registers\[26\]\[12\] net787 vssd1 vssd1 vccd1 vccd1 _02879_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1480_A a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13520__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06539_ cpu.f0.num\[12\] _01805_ _01812_ cpu.f0.i\[20\] _01910_ vssd1 vssd1 vccd1
+ vccd1 _01928_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14646__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09327_ _04212_ _04282_ _04284_ net493 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__o31a_1
XANTENNA__08076__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10958__A2 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__X _02162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ _03496_ _03497_ _03498_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or4_1
X_09189_ net302 net437 _04399_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_75_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_81_clk_X clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11220_ net1931 net190 net406 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10553__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__Q cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net2219 net195 net415 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
X_10102_ _05352_ _05372_ _05361_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o21a_1
XANTENNA__14026__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ net2718 net209 net425 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_96_clk_X clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09733__C1 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ net125 _05305_ _05309_ net627 vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a211o_1
XANTENNA__12113__X _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__C _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13050__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11984_ net2008 _05822_ net314 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09422__X _04713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A2 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ clknet_leaf_13_clk _00836_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10935_ cpu.DM0.readdata\[31\] _04447_ net734 vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13654_ clknet_leaf_61_clk _00767_ net1348 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_34_clk_X clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ cpu.DM0.readdata\[11\] net738 net722 vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__o21a_1
X_12605_ cpu.LCD0.row_2\[7\] net1789 net1012 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__mux2_1
XANTENNA__06925__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08067__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13585_ clknet_leaf_77_clk _00698_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10797_ cpu.f0.data_adr\[24\] _05107_ net993 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__mux2_1
XANTENNA__09803__A3 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ _06304_ _06305_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__nor2_1
XANTENNA__07814__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_clk_X clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ cpu.f0.i\[5\] _06260_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_91_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ clknet_leaf_85_clk _01319_ net1272 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11418_ net2643 net207 net382 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ cpu.DM0.data_i\[7\] net532 _05849_ _01791_ _01780_ vssd1 vssd1 vccd1 vccd1
+ _06222_ sky130_fd_sc_hd__a311o_2
XANTENNA__07578__A1 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14137_ clknet_leaf_42_clk _01250_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11349_ cpu.RF0.registers\[10\]\[13\] net197 net390 vssd1 vssd1 vccd1 vccd1 _00773_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14068_ clknet_leaf_71_clk _01181_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ clknet_leaf_36_clk _00208_ net1263 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
X_06890_ net1072 net1070 net1067 net1065 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and4bb_1
XANTENNA__06669__A a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__B1 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__X _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06553__A2 cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A1 cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ cpu.RF0.registers\[12\]\[5\] net697 net643 cpu.RF0.registers\[3\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a22o_1
XANTENNA__06956__X _02247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13543__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ net1057 cpu.RF0.registers\[18\]\[6\] net772 vssd1 vssd1 vccd1 vccd1 _02802_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08491_ cpu.RF0.registers\[18\]\[7\] net681 net641 cpu.RF0.registers\[19\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09699__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ net1055 cpu.RF0.registers\[19\]\[1\] net824 vssd1 vssd1 vccd1 vccd1 _02733_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_18_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07373_ net1054 cpu.RF0.registers\[23\]\[2\] net819 vssd1 vssd1 vccd1 vccd1 _02664_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09255__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__B2 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13693__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _04380_ _04395_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ net1027 cpu.RF0.registers\[17\]\[31\] net804 vssd1 vssd1 vccd1 vccd1 _04334_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_A _05799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13617__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__X _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 cpu.RF0.registers\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14049__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07666__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold421 cpu.RF0.registers\[0\]\[14\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 cpu.RF0.registers\[27\]\[2\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 cpu.RF0.registers\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 cpu.RF0.registers\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 cpu.RF0.registers\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 cpu.RF0.registers\[19\]\[31\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 cpu.RF0.registers\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _01940_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
Xhold498 cpu.RF0.registers\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 net914 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ cpu.IM0.address_IM\[9\] _05219_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__xor2_2
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_5_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 net937 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_A _02037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net951 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14199__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net961 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09226__Y _04517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ _05164_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__xor2_1
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_87_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 cpu.LCD0.row_1\[25\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
Xhold1121 _00331_ vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1132 cpu.RF0.registers\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ net1085 cpu.RF0.registers\[24\]\[19\] net870 vssd1 vssd1 vccd1 vccd1 _04118_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10876__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 cpu.LCD0.row_1\[75\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1154 _01618_ vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 cpu.RF0.registers\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 cpu.LCD0.row_1\[78\] vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 cpu.K0.count\[1\] vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _03669_ _04048_ _04046_ _04043_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_64_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 cpu.RF0.registers\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_07709_ net1037 cpu.RF0.registers\[31\]\[17\] net826 vssd1 vssd1 vccd1 vccd1 _03000_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08297__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08689_ cpu.RF0.registers\[7\]\[1\] net653 _03968_ _03970_ _03971_ vssd1 vssd1 vccd1
+ vccd1 _03980_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11424__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10720_ a1.ADR_I\[1\] net559 net537 _05690_ vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a22o_1
XANTENNA__12910__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07203__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__Q cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ net2705 cpu.LCD0.row_1\[65\] net906 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XANTENNA__09246__A1 _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12250__B1 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ _05678_ cpu.LCD0.row_1\[3\] net896 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
XANTENNA__09797__A2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13370_ clknet_leaf_93_clk _00483_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12321_ net1660 _05948_ _06199_ net1341 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12108__X _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__X _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ cpu.LCD0.row_1\[69\] _06001_ _06036_ cpu.LCD0.row_1\[21\] _06147_ vssd1 vssd1
+ vccd1 vccd1 _06148_ sky130_fd_sc_hd__a221o_1
XANTENNA__09403__D1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12553__B2 _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net2478 net236 net408 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12183_ _06064_ _06066_ _06068_ _06081_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__or4_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ cpu.RF0.registers\[3\]\[31\] net128 net418 vssd1 vssd1 vccd1 vccd1 _00567_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06783__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ net1848 net140 net428 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10016_ cpu.IM0.address_IM\[15\] _05284_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ net2436 net241 net316 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__mux2_1
XANTENNA__08288__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11334__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ clknet_leaf_102_clk _00819_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ net2133 net162 net432 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11898_ net1724 net253 net323 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13637_ clknet_leaf_8_clk _00750_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10849_ _05199_ _05782_ net721 vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__mux2_4
XANTENNA__12241__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13568_ clknet_leaf_3_clk _00681_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12519_ _01817_ _06293_ net260 vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06671__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13499_ clknet_leaf_12_clk _00612_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08460__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07486__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13096__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14341__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 net211 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _05790_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13909__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ net1093 cpu.RF0.registers\[28\]\[28\] net868 vssd1 vssd1 vccd1 vccd1 _03282_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11509__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _05019_ _05020_ net456 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__mux2_1
X_06942_ net954 cpu.RF0.registers\[14\]\[26\] net761 vssd1 vssd1 vccd1 vccd1 _02233_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10858__A1 _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14389__Q cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ _02866_ _03766_ _04840_ _03729_ _02545_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__o32a_1
X_06873_ net1067 net1065 net1072 net1069 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__and4b_1
XFILLER_0_94_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ net1101 cpu.RF0.registers\[21\]\[3\] _02019_ vssd1 vssd1 vccd1 vccd1 _03903_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12933__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ net292 _04485_ _04606_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__nor3_1
X_08543_ _02122_ _02796_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout161_A _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06846__B net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__A2 _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08474_ cpu.RF0.registers\[0\]\[8\] net664 net550 vssd1 vssd1 vccd1 vccd1 _03765_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08119__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07023__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ cpu.RF0.registers\[0\]\[0\] net618 _02699_ _02715_ vssd1 vssd1 vccd1 vccd1
+ _02716_ sky130_fd_sc_hd__o22a_2
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__X _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_A _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12232__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ net1055 cpu.RF0.registers\[31\]\[2\] net828 vssd1 vssd1 vccd1 vccd1 _02647_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_45_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07287_ _02569_ _02570_ _02576_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__nor4_1
XANTENNA__10384__A cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13439__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1335_A net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ cpu.RF0.registers\[12\]\[31\] net696 _04314_ _04315_ _04316_ vssd1 vssd1
+ vccd1 vccd1 _04317_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07396__C net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 cpu.FetchedInstr\[10\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 cpu.RF0.registers\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08203__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1123_X net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 cpu.RF0.registers\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 cpu.RF0.registers\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13589__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 cpu.RF0.registers\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 cpu.RF0.registers\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _02002_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11419__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_2
X_09928_ cpu.IM0.address_IM\[7\] net933 _05212_ _05213_ vssd1 vssd1 vccd1 vccd1 _00030_
+ sky130_fd_sc_hd__a22o_1
Xfanout753 _05639_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_2
Xfanout764 _02183_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_6
XANTENNA__09164__A0 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_4
Xfanout786 net787 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
X_09859_ _01785_ _02644_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nor2_1
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
XANTENNA__08020__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ clknet_leaf_5_clk cpu.c0.next_count\[1\] net1145 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11821_ net1671 net154 net334 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06756__B net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ clknet_leaf_46_clk _01642_ net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09132__B _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ net2867 net181 net344 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14214__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ cpu.LCD0.row_1\[109\] cpu.LCD0.row_1\[117\] net899 vssd1 vssd1 vccd1 vccd1
+ _00333_ sky130_fd_sc_hd__mux2_1
X_14471_ clknet_leaf_33_clk _01581_ net1250 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10846__X _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ net2545 net189 net350 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XANTENNA__08690__A2 _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ clknet_leaf_1_clk _00535_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ net2695 net2555 net909 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
XANTENNA__12223__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13353_ clknet_leaf_18_clk _00466_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_10565_ net59 net919 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__and2_1
XANTENNA__10785__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14364__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ net2814 net114 cpu.K0.next_state vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13284_ clknet_leaf_20_clk cpu.RU0.next_FetchedInstr\[23\] net1169 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[23\] sky130_fd_sc_hd__dfrtp_1
X_10496_ net1532 net916 net751 a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 _00169_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ net1420 net555 _06131_ net1354 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__o211a_1
XANTENNA__11268__A_N cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12166_ cpu.LCD0.row_2\[58\] _06000_ _06033_ cpu.LCD0.row_2\[74\] vssd1 vssd1 vccd1
+ vccd1 _06065_ sky130_fd_sc_hd__a22o_1
XANTENNA__11329__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ net1979 net193 net420 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__mux2_1
XANTENNA__12956__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _05995_ _05996_ net557 vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__and3_4
XANTENNA__09155__B1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ net2017 net209 net426 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__mux2_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08902__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12301__X _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ clknet_leaf_35_clk _00188_ net1258 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06666__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11999__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ net1391 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_28_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08681__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ cpu.RF0.registers\[14\]\[10\] net576 _02484_ _02488_ _02491_ vssd1 vssd1
+ vccd1 vccd1 _02501_ sky130_fd_sc_hd__a2111o_1
X_08190_ net939 cpu.RF0.registers\[3\]\[21\] net835 vssd1 vssd1 vccd1 vccd1 _03481_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08969__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ _02423_ _02424_ _02426_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__or4_2
XANTENNA__12765__B2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08433__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07072_ net974 cpu.RF0.registers\[4\]\[18\] net782 vssd1 vssd1 vccd1 vccd1 _02363_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12517__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13731__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09933__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11239__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ cpu.RF0.registers\[20\]\[29\] net709 _03262_ _03263_ _03264_ vssd1 vssd1
+ vccd1 vccd1 _03265_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14068__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13881__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09713_ _04360_ _04997_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a21oi_1
X_06925_ net1026 cpu.RF0.registers\[21\]\[26\] net795 vssd1 vssd1 vccd1 vccd1 _02216_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout376_A _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _02982_ _04159_ _04934_ _04933_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a31o_1
X_06856_ net1071 net1066 net1068 net1073 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06857__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13111__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07172__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14237__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ _03932_ _04399_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__or2_1
XANTENNA__09449__A1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06787_ cpu.RF0.registers\[27\]\[30\] net711 net646 cpu.RF0.registers\[21\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a22o_1
X_08526_ net1103 cpu.RF0.registers\[17\]\[6\] net885 vssd1 vssd1 vccd1 vccd1 _03817_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10059__A2 _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__B1 cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ net1095 cpu.RF0.registers\[21\]\[8\] net865 vssd1 vssd1 vccd1 vccd1 _03748_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13261__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14387__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11702__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ _02686_ _02690_ _02694_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08388_ net941 cpu.RF0.registers\[14\]\[10\] net838 vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10826__B cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12756__B2 cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07339_ net1064 cpu.RF0.registers\[26\]\[3\] net789 vssd1 vssd1 vccd1 vccd1 _02630_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_34_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08424__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07975__X _03266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ cpu.f0.i\[26\] _05579_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09619__A2_N _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ net1076 cpu.RF0.registers\[17\]\[31\] net882 vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__and3_1
X_10281_ cpu.f0.i\[15\] cpu.f0.i\[16\] _05518_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__and3_2
XANTENNA__12979__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ net1894 net177 net312 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__Q cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _02087_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
Xfanout561 _05686_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 _02189_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_8
Xfanout583 _02175_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_8
X_13971_ clknet_leaf_69_clk _01084_ net1326 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__A1 _04710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _02160_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_8
X_12922_ clknet_leaf_26_clk _00111_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12121__X _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07215__X _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ clknet_leaf_23_clk _00072_ net1194 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06910__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13604__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ net2031 net229 net337 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06917__D net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12784_ net1414 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14523_ clknet_leaf_61_clk net1585 net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_11735_ net1690 net247 net343 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08663__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11612__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07598__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14454_ clknet_leaf_25_clk _01564_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10470__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11666_ net1769 net238 net353 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XANTENNA__07871__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__A1 cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13754__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14492__Q cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06933__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13405_ clknet_leaf_88_clk _00518_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net2277 net2052 net904 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
X_14385_ clknet_leaf_24_clk _01496_ net1205 vssd1 vssd1 vccd1 vccd1 cpu.CU0.funct3\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11597_ net2710 net139 net362 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
X_13336_ clknet_leaf_18_clk _00449_ net1198 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10548_ net1133 net1792 net913 _05661_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__a31o_1
XANTENNA__06977__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13267_ clknet_leaf_34_clk cpu.RU0.next_FetchedInstr\[6\] net1247 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10479_ net1458 net922 net747 a1.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a22o_1
XANTENNA__08179__A1 cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ cpu.LCD0.row_2\[52\] _06011_ _06018_ cpu.LCD0.row_2\[100\] vssd1 vssd1 vccd1
+ vccd1 _06115_ sky130_fd_sc_hd__a22o_1
XANTENNA__09318__A _03119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A2 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ clknet_leaf_78_clk _00378_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11059__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12149_ _05981_ net744 net557 vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__and3_1
XANTENNA__14161__RESET_B net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13134__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__X _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10898__S net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06710_ _01999_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__and2_2
X_07690_ cpu.RF0.registers\[0\]\[16\] net617 _02976_ _02980_ vssd1 vssd1 vccd1 vccd1
+ _02981_ sky130_fd_sc_hd__o22a_2
XANTENNA__06677__A a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ a1.CPU_DAT_O\[9\] net895 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[9\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__13284__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _04521_ _04624_ _04650_ net470 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a22oi_2
X_06572_ cpu.c0.count\[1\] cpu.c0.count\[3\] cpu.c0.count\[2\] vssd1 vssd1 vccd1 vccd1
+ _01952_ sky130_fd_sc_hd__and3_1
X_08311_ net941 cpu.RF0.registers\[10\]\[12\] net861 vssd1 vssd1 vccd1 vccd1 _03602_
+ sky130_fd_sc_hd__and3_1
X_09291_ net470 _04374_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07004__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10997__A0 cpu.f0.write_data\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11522__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_13 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08242_ cpu.RF0.registers\[0\]\[14\] net664 net549 vssd1 vssd1 vccd1 vccd1 _03533_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_24 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_46 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__A1 cpu.f0.write_data\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__C net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08173_ net949 cpu.RF0.registers\[5\]\[20\] net865 vssd1 vssd1 vccd1 vccd1 _03464_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10749__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08406__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07124_ net969 cpu.RF0.registers\[2\]\[15\] net771 vssd1 vssd1 vccd1 vccd1 _02415_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06968__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ _02335_ _02336_ _02337_ _02345_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1033_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09906__A2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07674__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1200_A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ net1098 cpu.RF0.registers\[26\]\[29\] net861 vssd1 vssd1 vccd1 vccd1 _03248_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ cpu.RF0.registers\[26\]\[27\] net599 _02158_ _02178_ _02130_ vssd1 vssd1
+ vccd1 vccd1 _02199_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13627__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ cpu.RF0.registers\[23\]\[29\] net613 _02151_ cpu.RF0.registers\[29\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07145__A2 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09627_ _03145_ net446 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__xnor2_1
X_06839_ net1038 cpu.RF0.registers\[31\]\[27\] net827 vssd1 vssd1 vccd1 vccd1 _02130_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout925_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ _02865_ _03766_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08509_ _02582_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _04416_ _04423_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ net2050 net172 net373 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09410__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12825__Q cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13007__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ net2662 net205 net378 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
Xwire258 _05129_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_1
X_10402_ cpu.f0.i\[13\] net268 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nand2_1
X_14170_ clknet_leaf_94_clk _01283_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10204__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ net2811 net197 net386 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__mux2_1
X_13121_ clknet_leaf_47_clk _00301_ net1355 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[85\]
+ sky130_fd_sc_hd__dfstp_1
X_10333_ net1461 net724 _05479_ _05570_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13157__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ clknet_leaf_49_clk net2458 net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10264_ cpu.f0.i\[7\] cpu.f0.i\[13\] _05503_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__and3_1
XANTENNA__07584__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14402__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ net2380 net227 net313 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1301 net1313 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
Xfanout1312 net1313 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10912__A0 cpu.DM0.readdata\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ cpu.IM0.address_IM\[30\] _03232_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1323 net1326 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__clkbuf_4
Xfanout1334 net1335 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__buf_2
XANTENNA__07384__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1345 net1346 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1356 net1363 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__clkbuf_2
Xfanout1367 net1385 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__buf_2
Xfanout1378 net1384 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__clkbuf_4
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_4
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11607__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ clknet_leaf_10_clk _01067_ net1222 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14552__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07136__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ clknet_leaf_26_clk _00094_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06928__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13885_ clknet_leaf_67_clk _00998_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ clknet_leaf_33_clk _00055_ net1245 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08097__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ cpu.f0.write_data\[25\] net498 net279 cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1
+ _01746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A2 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ clknet_leaf_51_clk _01608_ net1377 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11718_ net1843 net172 net349 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ cpu.LCD0.row_2\[100\] cpu.LCD0.row_2\[92\] net1004 vssd1 vssd1 vccd1 vccd1
+ _01691_ sky130_fd_sc_hd__mux2_1
XANTENNA__07759__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14437_ clknet_leaf_15_clk net1122 net1243 vssd1 vssd1 vccd1 vccd1 cpu.IM0.pc_enable
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11649_ net2822 net207 net354 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12196__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14368_ clknet_leaf_57_clk _01481_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06960__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold806 cpu.RF0.registers\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold817 cpu.RF0.registers\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold828 _01637_ vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_18_clk cpu.RU0.next_FetchedData\[26\] net1192 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold839 cpu.RF0.registers\[23\]\[10\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
X_14299_ clknet_leaf_13_clk _01412_ net1241 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14082__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08860_ cpu.RF0.registers\[9\]\[16\] net699 net691 cpu.RF0.registers\[10\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1506 cpu.RF0.registers\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net2912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07791__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ net1032 cpu.RF0.registers\[21\]\[22\] net796 vssd1 vssd1 vccd1 vccd1 _03102_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1517 cpu.RF0.registers\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net2923 sky130_fd_sc_hd__dlygate4sd3_1
X_08791_ cpu.RF0.registers\[6\]\[18\] net676 _04057_ _04062_ _04067_ vssd1 vssd1 vccd1
+ vccd1 _04082_ sky130_fd_sc_hd__a2111o_1
Xhold1528 cpu.LCD0.row_1\[54\] vssd1 vssd1 vccd1 vccd1 net2934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11517__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07742_ cpu.RF0.registers\[22\]\[20\] net604 net600 cpu.RF0.registers\[26\]\[20\]
+ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07127__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06838__C net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14397__Q cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07673_ net1024 cpu.RF0.registers\[31\]\[16\] net825 vssd1 vssd1 vccd1 vccd1 _02964_
+ sky130_fd_sc_hd__and3_1
X_09412_ _03172_ net435 _04701_ net294 net289 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__o221a_1
X_06624_ _01970_ _01990_ _01991_ _01971_ _01986_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09511__A _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _04456_ _04500_ net470 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__mux2_1
X_06555_ cpu.f0.state\[8\] _01871_ _01941_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout241_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07835__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _04371_ _04564_ _04563_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07669__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06486_ cpu.FetchedInstr\[17\] cpu.FetchedInstr\[16\] cpu.FetchedInstr\[19\] cpu.FetchedInstr\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08225_ cpu.RF0.registers\[15\]\[14\] net683 net648 cpu.RF0.registers\[25\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1150_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__A2 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08156_ _03443_ _03444_ _03445_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07107_ cpu.RF0.registers\[7\]\[14\] net595 net591 cpu.RF0.registers\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10392__A cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ net1082 cpu.RF0.registers\[30\]\[22\] net837 vssd1 vssd1 vccd1 vccd1 _03378_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07038_ net1041 cpu.RF0.registers\[27\]\[19\] net776 vssd1 vssd1 vccd1 vccd1 _02329_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06869__X _02160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09245__X _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10370__A1 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _04243_ _04245_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__and2_1
XANTENNA__11427__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _02579_ net515 vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10122__A1 cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08866__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ clknet_leaf_6_clk _00783_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ net723 _05294_ _05805_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a22o_2
XFILLER_0_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ net2465 net2631 net1004 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
XANTENNA__08963__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__B2 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ cpu.f0.state\[8\] _01872_ cpu.f0.next_write_i _06319_ vssd1 vssd1 vccd1 vccd1
+ _06320_ sky130_fd_sc_hd__a211o_4
XANTENNA__09140__B _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07579__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11503_ net1742 net249 net371 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__mux2_1
X_12483_ net263 _06271_ _06272_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__and3_1
XANTENNA__12178__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14222_ clknet_leaf_2_clk _01335_ net1154 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11434_ _05766_ net503 _05910_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ clknet_leaf_105_clk _01266_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08251__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_100_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11365_ net2639 net142 net391 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__mux2_1
X_13104_ clknet_leaf_49_clk _00284_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[68\]
+ sky130_fd_sc_hd__dfstp_1
X_10316_ cpu.f0.i\[21\] _05549_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14084_ clknet_leaf_96_clk _01197_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11296_ net2069 net157 net398 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ clknet_leaf_31_clk _00013_ net1205 vssd1 vssd1 vccd1 vccd1 cpu.DM0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ cpu.f0.i\[11\] _05491_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and2_1
XANTENNA__11689__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_2
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_clk_X clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__A1 cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1153 net1154 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ cpu.IM0.address_IM\[28\] cpu.IM0.address_IM\[27\] _05422_ vssd1 vssd1 vccd1
+ vccd1 _05443_ sky130_fd_sc_hd__and3_2
XFILLER_0_101_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11337__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_4
Xfanout1175 net1191 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_59_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1186 net1191 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_2
XANTENNA__07109__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ clknet_leaf_77_clk _01050_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09034__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13868_ clknet_leaf_74_clk _00981_ net1324 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ clknet_leaf_16_clk _00038_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13799_ clknet_leaf_81_clk _00912_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06674__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11072__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07489__C net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13322__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14448__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08490__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11800__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ _03150_ _03172_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06690__A a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__A3 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 cpu.RF0.registers\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 cpu.RF0.registers\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold625 cpu.RF0.registers\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13472__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14598__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold636 cpu.RF0.registers\[22\]\[23\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _00255_ vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 cpu.RF0.registers\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire843_A _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ _05242_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__nor2_1
Xhold669 cpu.RF0.registers\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload26_A clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ _04055_ _04056_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09892_ net127 _05180_ _05177_ net631 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a211o_1
XANTENNA__09742__A0 _04396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07348__A2 _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net1074 cpu.RF0.registers\[29\]\[16\] net848 vssd1 vssd1 vccd1 vccd1 _04134_
+ sky130_fd_sc_hd__and3_1
Xhold1303 cpu.RF0.registers\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07952__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1314 cpu.LCD0.row_1\[80\] vssd1 vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11247__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1325 cpu.RF0.registers\[0\]\[28\] vssd1 vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1336 cpu.RF0.registers\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08774_ net948 cpu.RF0.registers\[15\]\[18\] net858 vssd1 vssd1 vccd1 vccd1 _04065_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1347 cpu.RF0.registers\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 cpu.RF0.registers\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1369 cpu.RF0.registers\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07725_ cpu.RF0.registers\[10\]\[17\] net569 _02988_ _02991_ _02993_ vssd1 vssd1
+ vccd1 vccd1 _03016_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_36_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10104__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1198_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ net1115 _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06865__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__B cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06607_ _01972_ _01755_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ net1046 cpu.RF0.registers\[29\]\[12\] net792 vssd1 vssd1 vccd1 vccd1 _02878_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1365_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ net512 _04554_ _04602_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o31a_2
XFILLER_0_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06538_ cpu.f0.num\[2\] _01792_ _01802_ cpu.f0.i\[11\] _01916_ vssd1 vssd1 vccd1
+ vccd1 _01927_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ net305 _04523_ _04527_ _04547_ _04542_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__o221a_1
X_06469_ cpu.DM0.enable _01849_ cpu.DM0.state\[0\] vssd1 vssd1 vccd1 vccd1 _01865_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11710__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08208_ cpu.RF0.registers\[16\]\[21\] net636 _03480_ _03482_ _03484_ vssd1 vssd1
+ vccd1 vccd1 _03499_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ net302 net437 _04399_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09025__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout992_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08233__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ cpu.RF0.registers\[14\]\[23\] net650 _03427_ _03428_ _03429_ vssd1 vssd1
+ vccd1 vccd1 _03430_ sky130_fd_sc_hd__a2111o_1
X_11150_ net2176 net197 net414 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13965__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ cpu.IM0.address_IM\[20\] _03042_ _03078_ cpu.IM0.address_IM\[21\] vssd1 vssd1
+ vccd1 vccd1 _05372_ sky130_fd_sc_hd__a22o_1
X_11081_ net2417 net203 net422 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ net715 net132 _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and3_1
XANTENNA__06547__B1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11157__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__B net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__X _05783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__C1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ net2735 net182 net317 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__mux2_1
X_13722_ clknet_leaf_90_clk _00835_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10934_ net1886 net137 net430 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__mux2_1
XANTENNA__06775__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13345__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13653_ clknet_leaf_73_clk _00766_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10865_ _01852_ _04792_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or2_1
XANTENNA__10297__A cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ cpu.LCD0.row_2\[6\] net1645 net1012 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__mux2_1
XANTENNA__12399__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13584_ clknet_leaf_74_clk _00697_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10796_ a1.ADR_I\[23\] net558 net536 _05744_ vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12535_ _01821_ _06303_ net260 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13495__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11620__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ _06260_ _06261_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nor2_1
XANTENNA__09016__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06941__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ clknet_leaf_67_clk _01318_ net1294 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11417_ net2888 net173 net385 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08224__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ net1546 cpu.DM0.data_i\[7\] cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1 _01523_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07578__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14136_ clknet_leaf_7_clk _01249_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ net1781 net210 net393 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XANTENNA__10582__A1 cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_68_clk _01180_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11279_ net2454 net217 net398 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__mux2_1
X_13018_ clknet_leaf_34_clk _00207_ net1252 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10334__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06669__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11067__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__X _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07510_ net978 cpu.RF0.registers\[9\]\[6\] net760 vssd1 vssd1 vccd1 vccd1 _02801_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ cpu.RF0.registers\[12\]\[7\] net697 net669 cpu.RF0.registers\[22\]\[7\] _03776_
+ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07441_ net1058 cpu.RF0.registers\[25\]\[1\] net760 vssd1 vssd1 vccd1 vccd1 _02732_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_18_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13838__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ net1054 cpu.RF0.registers\[17\]\[2\] net807 vssd1 vssd1 vccd1 vccd1 _02663_
+ sky130_fd_sc_hd__and3_1
X_09111_ _04380_ _04395_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__nor2_4
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11530__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ net954 cpu.RF0.registers\[13\]\[31\] net790 vssd1 vssd1 vccd1 vccd1 _04333_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_72_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12862__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06851__C net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13988__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07018__A1 cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 _00290_ vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 cpu.RF0.registers\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09412__C1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 cpu.RU0.state\[2\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _05796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07569__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 cpu.RF0.registers\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__B1 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold444 cpu.FetchedInstr\[21\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 cpu.RF0.registers\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 cpu.RF0.registers\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 a1.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net905 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
X_09944_ _05226_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__xnor2_1
Xhold488 cpu.RF0.registers\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13218__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_2
Xhold499 cpu.RF0.registers\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 _01859_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_2
XANTENNA__08778__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net951 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09236__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _05151_ _05156_ _05150_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a21o_1
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 cpu.RF0.registers\[16\]\[31\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net984 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _00249_ vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net983 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_2
Xhold1122 cpu.LCD0.row_1\[33\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net1085 cpu.RF0.registers\[18\]\[19\] net855 vssd1 vssd1 vccd1 vccd1 _04117_
+ sky130_fd_sc_hd__and3_1
Xhold1133 cpu.RF0.registers\[0\]\[7\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 cpu.RF0.registers\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 cpu.RF0.registers\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07741__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13368__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 cpu.RF0.registers\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _03668_ _04041_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2_1
Xhold1177 _00302_ vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14613__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 cpu.RF0.registers\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 cpu.LCD0.row_2\[78\] vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11705__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _02052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ net952 cpu.RF0.registers\[15\]\[17\] net825 vssd1 vssd1 vccd1 vccd1 _02999_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08688_ cpu.RF0.registers\[4\]\[1\] net679 net647 cpu.RF0.registers\[21\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ cpu.RF0.registers\[2\]\[13\] net584 _02909_ _02911_ _02924_ vssd1 vssd1 vccd1
+ vccd1 _02930_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ net2370 cpu.LCD0.row_1\[64\] net909 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XANTENNA__06882__X _02173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08018__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _04589_ _04592_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10581_ cpu.f0.write_data\[3\] _02641_ net996 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08454__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11440__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12320_ _05951_ _05956_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__or2_1
XANTENNA__08315__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12833__Q cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ cpu.LCD0.row_2\[93\] _05983_ _06021_ cpu.LCD0.row_1\[93\] vssd1 vssd1 vccd1
+ vccd1 _06147_ sky130_fd_sc_hd__a22o_1
XANTENNA__08206__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ net504 _05912_ _05915_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__and3_4
X_12182_ cpu.LCD0.row_1\[122\] _06014_ _06070_ _06080_ net556 vssd1 vssd1 vccd1 vccd1
+ _06081_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10564__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net2698 net137 net418 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XANTENNA__14143__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__X _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net2419 net144 net428 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XANTENNA__07592__C _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10015_ _05291_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08985__A _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14293__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11615__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ net1625 net247 net316 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14495__Q cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06936__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ clknet_leaf_104_clk _00818_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10917_ net723 _05413_ _05830_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_15_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11897_ net1753 net238 net324 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13636_ clknet_leaf_99_clk _00749_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10848_ cpu.DM0.readdata\[6\] _04896_ net739 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12885__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ clknet_leaf_2_clk _00680_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08445__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ net991 _04683_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11350__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12518_ net1018 cpu.f0.i\[24\] _06291_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07767__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13498_ clknet_leaf_96_clk _00611_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12449_ net1129 _06248_ net309 vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14119_ clknet_leaf_81_clk _01232_ net1291 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_07990_ net945 cpu.RF0.registers\[2\]\[28\] net854 vssd1 vssd1 vccd1 vccd1 _03281_
+ sky130_fd_sc_hd__and3_1
Xfanout209 net211 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07971__A2 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ net1029 cpu.RF0.registers\[29\]\[26\] net790 vssd1 vssd1 vccd1 vccd1 _02232_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10307__A1 _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14636__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ _04815_ _04816_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__and2b_1
X_06872_ net1038 cpu.RF0.registers\[21\]\[27\] net796 vssd1 vssd1 vccd1 vccd1 _02163_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _03899_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__and2_1
X_09591_ _03870_ _04035_ _04036_ _03836_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07007__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ cpu.IM0.address_IM\[6\] net553 _03831_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_
+ sky130_fd_sc_hd__a22o_2
XANTENNA__12210__A _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload93_A clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06846__C net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _03740_ _03747_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout154_A _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _02703_ _02706_ _02710_ _02714_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14016__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_clk_X clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07355_ net976 cpu.RF0.registers\[1\]\[2\] net807 vssd1 vssd1 vccd1 vccd1 _02646_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout321_A _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11260__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout419_A _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ cpu.RF0.registers\[20\]\[7\] net594 _02564_ _02567_ _02568_ vssd1 vssd1 vccd1
+ vccd1 _02577_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10384__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__A1 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09025_ cpu.RF0.registers\[11\]\[31\] net690 net687 cpu.RF0.registers\[31\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14166__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1230_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1328_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 cpu.RF0.registers\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold241 cpu.RF0.registers\[22\]\[18\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10546__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_A _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 cpu.RF0.registers\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 cpu.RF0.registers\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 cpu.LCD0.row_1\[122\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 cpu.RF0.registers\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 cpu.RF0.registers\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _02011_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_33_clk_X clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_4
XANTENNA__13190__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_2
XANTENNA__07962__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ net631 _04880_ net933 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a21oi_1
Xfanout743 _05985_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_2
Xfanout754 _05638_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net768 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09164__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout776 net779 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
X_09858_ net716 net132 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout787 net789 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
XANTENNA__07175__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout798 _02147_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_8
X_08809_ net938 cpu.RF0.registers\[13\]\[19\] net849 vssd1 vssd1 vccd1 vccd1 _04100_
+ sky130_fd_sc_hd__and3_1
X_09789_ _02410_ net435 net289 _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_48_clk_X clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11435__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11820_ net2604 net165 net334 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__mux2_1
XANTENNA__09467__A2 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12828__Q cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11751_ net1543 net171 net342 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__mux2_1
XANTENNA__12471__A1 cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
X_10702_ cpu.LCD0.row_1\[108\] cpu.LCD0.row_1\[116\] net903 vssd1 vssd1 vccd1 vccd1
+ _00332_ sky130_fd_sc_hd__mux2_1
X_14470_ clknet_leaf_34_clk _01580_ net1251 vssd1 vssd1 vccd1 vccd1 cpu.SR1.char_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11682_ net1783 net206 net350 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13421_ clknet_leaf_103_clk _00534_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ net2595 net2441 net905 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
XANTENNA__11026__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_106_clk_X clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11170__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06772__B _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14509__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ clknet_leaf_97_clk _00465_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ net1134 a1.ADR_I\[26\] net914 _05669_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__a31o_1
XANTENNA__07587__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10785__B2 _05736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net2801 net113 cpu.K0.next_state vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__mux2_1
X_13283_ clknet_leaf_20_clk cpu.RU0.next_FetchedInstr\[22\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[22\] sky130_fd_sc_hd__dfrtp_1
X_10495_ net1496 net916 net751 a1.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 _00168_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12790__A cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ _06111_ _06123_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__or3_1
XANTENNA__09927__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13533__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ cpu.LCD0.row_2\[10\] _05998_ _06012_ cpu.LCD0.row_2\[106\] _06063_ vssd1
+ vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11116_ net1749 net199 net419 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__mux2_1
X_12096_ _01773_ cpu.LCD0.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and2_1
XANTENNA__09155__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ net2051 net201 net427 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__mux2_1
XANTENNA__13683__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11345__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12998_ clknet_leaf_28_clk _00187_ net1201 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XANTENNA__14039__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07124__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__A1 cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ net1899 net172 net319 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08130__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14668_ net1390 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08881__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ clknet_leaf_69_clk _00732_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11017__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13063__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14189__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14599_ clknet_leaf_55_clk net2267 net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11080__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06682__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10225__B1 _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _02427_ _02428_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10776__A1 _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07071_ net1063 cpu.RF0.registers\[20\]\[18\] net782 vssd1 vssd1 vccd1 vccd1 _02362_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12900__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ cpu.RF0.registers\[8\]\[29\] net707 net701 cpu.RF0.registers\[9\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a22o_1
X_09712_ _04380_ _04405_ _04990_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__or4bb_1
XANTENNA__08121__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06924_ net1026 cpu.RF0.registers\[30\]\[26\] net761 vssd1 vssd1 vccd1 vccd1 _02215_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12150__B1 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _03019_ net439 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06855_ net1059 net802 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07960__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06857__B net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _04038_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__xor2_2
XANTENNA__12813__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06786_ cpu.RF0.registers\[5\]\[30\] net702 net640 cpu.RF0.registers\[19\]\[30\]
+ _02048_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09449__A2 _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net949 cpu.RF0.registers\[14\]\[6\] net840 vssd1 vssd1 vccd1 vccd1 _03816_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12453__A1 cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__C1 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_60_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1278_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _03744_ _03745_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07407_ cpu.RF0.registers\[9\]\[0\] net574 _02695_ _02696_ _02697_ vssd1 vssd1 vccd1
+ vccd1 _02698_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11008__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ cpu.RF0.registers\[5\]\[10\] net703 net669 cpu.RF0.registers\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ net974 cpu.RF0.registers\[7\]\[3\] net818 vssd1 vssd1 vccd1 vccd1 _02629_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10767__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13556__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__B2 cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07200__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ net980 cpu.RF0.registers\[2\]\[7\] net772 vssd1 vssd1 vccd1 vccd1 _02560_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09008_ net934 cpu.RF0.registers\[6\]\[31\] net851 vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__and3_1
X_10280_ cpu.f0.i\[15\] _05518_ cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A1 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_4
Xfanout562 _05641_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
Xfanout573 _02187_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_8
X_13970_ clknet_leaf_60_clk _01083_ net1344 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout584 _02173_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_13_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08966__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_25_clk _00110_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08896__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11165__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12852_ clknet_leaf_39_clk _00071_ net1254 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net2521 net233 net337 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ net1554 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13086__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14522_ clknet_leaf_51_clk _01624_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_11734_ net1895 net249 net344 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14453_ clknet_leaf_24_clk _01563_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07871__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ net505 _05906_ _05915_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__and3_4
XANTENNA__10207__B1 cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10616_ net2762 net2654 net907 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13404_ clknet_leaf_11_clk _00517_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07608__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14384_ clknet_leaf_23_clk _01495_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_11596_ net1673 net141 net364 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13335_ clknet_leaf_42_clk _00448_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ net49 net920 vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__and2_1
XANTENNA__08820__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[5\] net1246 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[5\] sky130_fd_sc_hd__dfrtp_1
X_10478_ net72 net915 _01861_ vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__o21a_1
X_12217_ cpu.LCD0.row_2\[84\] _05990_ _06003_ cpu.LCD0.row_2\[20\] _06113_ vssd1 vssd1
+ vccd1 vccd1 _06114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13197_ clknet_leaf_74_clk _00377_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09318__B _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ cpu.LCD0.row_1\[81\] _05986_ _06007_ cpu.LCD0.row_2\[113\] _06047_ vssd1
+ vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a221o_1
XANTENNA__09037__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12079_ cpu.LCD0.nextState\[5\] cpu.LCD0.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05980_
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06958__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08876__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08887__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06677__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13429__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06640_ a1.CPU_DAT_O\[8\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[8\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06571_ cpu.DM0.dhit _01791_ _01947_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08639__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__C1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08310_ net442 _03597_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__xor2_1
XANTENNA__08103__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07789__A _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__B2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ net470 _04572_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nand2_1
XANTENNA__06693__A a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13579__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07311__B1 _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ _03518_ _03520_ _03527_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_14 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__B1 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_47 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ cpu.RF0.registers\[9\]\[20\] net701 _03460_ _03461_ _03462_ vssd1 vssd1 vccd1
+ vccd1 _03463_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06843__D net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13299__Q cpu.DM0.data_i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__A2 _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__B2 cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ cpu.RF0.registers\[10\]\[15\] net570 _02191_ cpu.RF0.registers\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07054_ cpu.RF0.registers\[1\]\[19\] net588 net568 cpu.RF0.registers\[25\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a22o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__07955__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08413__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__12931__Q a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout486_A _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ net947 cpu.RF0.registers\[15\]\[29\] net858 vssd1 vssd1 vccd1 vccd1 _03247_
+ sky130_fd_sc_hd__and3_1
X_06907_ cpu.RF0.registers\[22\]\[27\] net604 _02152_ _02166_ _02142_ vssd1 vssd1
+ vccd1 vccd1 _02198_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07887_ cpu.RF0.registers\[8\]\[29\] net612 net602 cpu.RF0.registers\[5\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14354__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06838_ net1073 net1070 net1068 net1066 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__and4_4
X_09626_ _03146_ net446 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__nand2_1
X_09557_ _02865_ _03766_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nor2_1
X_06769_ net1080 cpu.RF0.registers\[25\]\[30\] net862 vssd1 vssd1 vccd1 vccd1 _02060_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout820_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11713__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08508_ _02796_ _02830_ _02122_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07699__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09488_ _04583_ _04778_ net302 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07302__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ _02832_ _02866_ net491 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11021__B1_N net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12946__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ net1901 net174 net379 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10401_ _01804_ net269 _05618_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08026__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11381_ net1702 net208 net389 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__mux2_1
XANTENNA__09070__A3 _03233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13120_ clknet_leaf_48_clk _00300_ net1361 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_10332_ net527 _05566_ _05569_ net307 vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08148__B1_N net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07081__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ clknet_leaf_47_clk _00231_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10263_ _05509_ _05510_ net309 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__or3b_1
XANTENNA__09138__B _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net2880 net231 net313 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__mux2_1
Xfanout1302 net1313 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
X_10194_ cpu.IM0.address_IM\[29\] net933 _05456_ _05457_ vssd1 vssd1 vccd1 vccd1 _00052_
+ sky130_fd_sc_hd__a22o_1
Xfanout1313 net1386 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10912__A1 _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1324 net1326 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1335 net1336 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__clkbuf_2
Xfanout1346 net1364 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1357 net1358 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12132__X _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout370 net373 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_6
Xfanout1368 net1371 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__buf_2
Xfanout1379 net1384 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__clkbuf_2
Xfanout381 _05926_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_8
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13953_ clknet_leaf_60_clk _01066_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ clknet_leaf_26_clk _00093_ net1181 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ clknet_leaf_15_clk _00997_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12835_ clknet_leaf_16_clk _00054_ net1243 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13721__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12719__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11623__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12766_ cpu.f0.write_data\[24\] net497 net279 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1
+ _01745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10747__B _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10979__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06944__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ clknet_leaf_49_clk net2195 net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11717_ net2005 net185 net348 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__mux2_1
XANTENNA__10239__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ net2306 cpu.LCD0.row_2\[91\] net998 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11648_ net2206 net174 net357 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__mux2_1
X_14436_ clknet_leaf_16_clk net2039 net1199 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11579_ net2598 net211 net362 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__mux2_1
X_14367_ clknet_leaf_57_clk _01480_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10600__A0 cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold807 cpu.RF0.registers\[28\]\[26\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold818 cpu.RF0.registers\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[25\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[25\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09329__A _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13101__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 cpu.LCD0.row_1\[106\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_93_clk _01411_ net1241 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14227__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13249_ clknet_leaf_35_clk _00429_ net1260 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10903__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__Y _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ net1031 cpu.RF0.registers\[29\]\[22\] net791 vssd1 vssd1 vccd1 vccd1 _03101_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13251__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14377__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1507 cpu.RF0.registers\[4\]\[23\] vssd1 vssd1 vccd1 vccd1 net2913 sky130_fd_sc_hd__dlygate4sd3_1
X_08790_ cpu.RF0.registers\[9\]\[18\] net700 net681 cpu.RF0.registers\[18\]\[18\]
+ _04070_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a221o_1
Xhold1518 cpu.RF0.registers\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net2924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06688__A a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1529 cpu.RF0.registers\[29\]\[2\] vssd1 vssd1 vccd1 vccd1 net2935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12819__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ cpu.RF0.registers\[8\]\[20\] net612 net593 cpu.RF0.registers\[21\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a22o_1
XANTENNA__08324__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ net953 cpu.RF0.registers\[3\]\[16\] net820 vssd1 vssd1 vccd1 vccd1 _02963_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06838__D net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ net298 _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__nand2_1
X_06623_ _01757_ _01984_ _01989_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12629__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12969__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ net449 _04511_ _04510_ _02758_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__o211ai_1
X_06554_ _01875_ _01886_ _01776_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08408__A _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07312__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__C net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ net484 _04383_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06485_ cpu.FetchedInstr\[21\] cpu.FetchedInstr\[20\] cpu.FetchedInstr\[23\] cpu.FetchedInstr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08224_ cpu.RF0.registers\[2\]\[14\] net655 net646 cpu.RF0.registers\[21\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ cpu.RF0.registers\[27\]\[20\] net712 net706 cpu.RF0.registers\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout401_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1143_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07106_ _02392_ _02394_ _02395_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__or4_1
X_08086_ net1080 cpu.RF0.registers\[19\]\[22\] net835 vssd1 vssd1 vccd1 vccd1 _03377_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10392__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ net1040 cpu.RF0.registers\[26\]\[19\] net789 vssd1 vssd1 vccd1 vccd1 _02328_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10960__X _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1310_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_A _02172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _04246_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13744__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ _03226_ _03228_ _03229_ _03199_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ net532 _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ net513 _04393_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ cpu.DM0.readdata\[15\] net735 net719 vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12620_ net2497 cpu.LCD0.row_2\[14\] net1006 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__mux2_1
XANTENNA__13894__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__A1 cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08318__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06764__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ _01780_ cpu.f0.state\[3\] net729 _06318_ vssd1 vssd1 vccd1 vccd1 _06319_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12836__Q cpu.f0.data_adr\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net2106 net256 net372 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__mux2_1
XANTENNA__10830__B1 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12482_ net541 net257 vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__nand2_1
XANTENNA__09028__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13124__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14221_ clknet_leaf_105_clk _01334_ net1156 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11433_ net1799 net131 net382 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12127__X _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ clknet_leaf_97_clk _01265_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07054__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ net2205 net146 net392 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08053__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ clknet_leaf_46_clk _00283_ net1356 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_10315_ net540 _05549_ cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13274__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14083_ clknet_leaf_78_clk _01196_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11295_ net1876 net161 net399 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ clknet_leaf_31_clk _00012_ net1205 vssd1 vssd1 vccd1 vccd1 cpu.DM0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10246_ _05496_ _05493_ net725 cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1 _00065_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_37_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1110 cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
XANTENNA__11618__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1121 cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_2
Xfanout1132 _01790_ vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_10177_ net718 net135 _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a21oi_1
Xfanout1143 net1211 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1154 net1167 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_2
XANTENNA__12549__A_N cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1176 net1180 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
Xfanout1187 net1191 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
X_13936_ clknet_leaf_74_clk _01049_ net1321 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10758__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ clknet_leaf_89_clk _00980_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11353__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ clknet_leaf_40_clk _00037_ net1243 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_6_clk _00911_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12749_ net1787 net498 net279 net1021 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09050__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10821__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07293__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ clknet_leaf_40_clk _01530_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06690__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold604 cpu.RF0.registers\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07045__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold615 cpu.RF0.registers\[17\]\[0\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold626 cpu.RF0.registers\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold637 cpu.RF0.registers\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold648 cpu.RF0.registers\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ cpu.IM0.address_IM\[9\] _05219_ cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1
+ vccd1 _05243_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10780__X _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold659 cpu.RF0.registers\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _04128_ _04165_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__or3_1
X_09891_ _05178_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nor2_1
XANTENNA__13767__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ net934 cpu.RF0.registers\[11\]\[16\] net880 vssd1 vssd1 vccd1 vccd1 _04133_
+ sky130_fd_sc_hd__and3_1
Xhold1304 cpu.RF0.registers\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 cpu.RF0.registers\[5\]\[6\] vssd1 vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 cpu.f0.num\[9\] vssd1 vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06849__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1337 cpu.LCD0.row_1\[49\] vssd1 vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ net1100 cpu.RF0.registers\[19\]\[18\] net836 vssd1 vssd1 vccd1 vccd1 _04064_
+ sky130_fd_sc_hd__and3_1
Xhold1348 cpu.RF0.registers\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 cpu.RF0.registers\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout184_A _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ cpu.RF0.registers\[28\]\[17\] net578 _02985_ _02992_ net621 vssd1 vssd1 vccd1
+ vccd1 _03015_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10104__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ _02832_ _02868_ _02944_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_81_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout351_A _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _01755_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__inv_2
XANTENNA__07313__Y _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ net968 cpu.RF0.registers\[12\]\[12\] net766 vssd1 vssd1 vccd1 vccd1 _02877_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13147__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _04496_ _04607_ _04613_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a211oi_2
X_06537_ cpu.f0.num\[18\] _01811_ _01816_ cpu.f0.i\[24\] _01917_ vssd1 vssd1 vccd1
+ vccd1 _01926_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1358_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10812__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ net278 _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nand2_1
X_06468_ _01788_ a1.READ_I a1.curr_state\[0\] net1135 a1.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _00009_ sky130_fd_sc_hd__a32o_1
XANTENNA__06881__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08207_ cpu.RF0.registers\[27\]\[21\] net711 net648 cpu.RF0.registers\[25\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13297__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ _04463_ _04477_ net484 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__mux2_1
X_06399_ net2906 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08138_ cpu.RF0.registers\[20\]\[23\] net710 net691 cpu.RF0.registers\[10\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout985_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ cpu.RF0.registers\[17\]\[25\] net694 _03348_ _03349_ _03354_ vssd1 vssd1
+ vccd1 vccd1 _03360_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1313_X net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10100_ _05369_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__and2b_1
X_11080_ net1764 net214 net424 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ _05306_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nor2_1
XANTENNA__09733__B2 _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07744__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11982_ net1707 net170 net314 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__mux2_1
X_13721_ clknet_leaf_92_clk _00834_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _05466_ _05842_ net719 vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06775__B net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10864_ net1728 net213 net432 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
X_13652_ clknet_leaf_71_clk _00765_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14072__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ cpu.LCD0.row_2\[5\] net1538 net1012 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ cpu.IM0.address_IM\[23\] net1013 net284 _05743_ vssd1 vssd1 vccd1 vccd1 _05744_
+ sky130_fd_sc_hd__a22o_1
X_13583_ clknet_leaf_82_clk _00696_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11901__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10803__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12534_ _01821_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10584__Y _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ cpu.f0.i\[4\] _06258_ net261 vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14204_ clknet_leaf_15_clk _01317_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11416_ net2104 net193 net385 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
X_12396_ net2278 cpu.DM0.data_i\[6\] net733 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11347_ net2049 net202 net392 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14135_ clknet_leaf_64_clk _01248_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_89_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11278_ net2800 net220 net400 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__mux2_1
X_14066_ clknet_leaf_60_clk _01179_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ clknet_leaf_29_clk _00206_ net1203 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09724__B2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ net1021 cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__nand2_1
XANTENNA__06538__B2 cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B1 _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13956__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 cpu.K0.state vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09045__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08884__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_106_clk _01032_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06685__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08160__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07440_ net977 cpu.RF0.registers\[3\]\[1\] net824 vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07371_ net976 cpu.RF0.registers\[4\]\[2\] net783 vssd1 vssd1 vccd1 vccd1 _02662_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ net437 _04399_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11811__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14565__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ net1025 cpu.RF0.registers\[22\]\[31\] net799 vssd1 vssd1 vccd1 vccd1 _04332_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07018__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 cpu.RF0.registers\[28\]\[6\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 cpu.RF0.registers\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 cpu.RF0.registers\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08124__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold434 cpu.RF0.registers\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold445 cpu.RF0.registers\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold456 cpu.RF0.registers\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 cpu.RF0.registers\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 cpu.RF0.registers\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ cpu.IM0.address_IM\[8\] _02833_ _05216_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a21o_1
Xhold489 cpu.RF0.registers\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout903 net905 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
Xfanout914 _01860_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout925 net929 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout399_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
X_09874_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__and2b_1
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_2
XANTENNA__11522__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout958 net960 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 cpu.RF0.registers\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 net984 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1106_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09804__X _05095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 cpu.RF0.registers\[22\]\[6\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net1084 cpu.RF0.registers\[26\]\[19\] net860 vssd1 vssd1 vccd1 vccd1 _04116_
+ sky130_fd_sc_hd__and3_1
Xhold1123 cpu.RF0.registers\[0\]\[17\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 cpu.RF0.registers\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 cpu.LCD0.row_2\[51\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 cpu.RF0.registers\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 cpu.RF0.registers\[0\]\[21\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _03735_ _03771_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__nor3_1
Xhold1178 cpu.RF0.registers\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 cpu.LCD0.row_1\[39\] vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ net959 cpu.RF0.registers\[11\]\[17\] net776 vssd1 vssd1 vccd1 vccd1 _02998_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout733_A cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08687_ cpu.RF0.registers\[28\]\[1\] net706 _02030_ cpu.RF0.registers\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07638_ cpu.RF0.registers\[21\]\[13\] net593 _02915_ _02917_ _02918_ vssd1 vssd1
+ vccd1 vccd1 _02929_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07569_ cpu.RF0.registers\[4\]\[8\] net587 _02845_ _02847_ _02853_ vssd1 vssd1 vccd1
+ vccd1 _02860_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07203__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09398__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _04414_ _04596_ _04598_ _04480_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a22oi_1
X_10580_ _05677_ cpu.LCD0.row_1\[2\] net901 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12250__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_clk_X clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13932__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _04417_ _04425_ net451 vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ cpu.LCD0.row_1\[109\] _06009_ _06019_ cpu.LCD0.row_1\[53\] _06145_ vssd1
+ vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07009__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11201_ net2890 net129 net410 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _06072_ _06074_ _06077_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__or4_1
XANTENNA__10861__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net2221 net142 net421 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
Xhold990 cpu.LCD0.row_2\[105\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ net1839 net151 net427 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
XANTENNA__09714__X _05005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _05278_ _05281_ _05276_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a21bo_1
XANTENNA__14438__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ net2935 net251 net317 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14588__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13704_ clknet_leaf_85_clk _00817_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10916_ cpu.DM0.readdata\[25\] net734 net719 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__o21a_1
X_14684_ net1406 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__07496__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B1 cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11896_ net506 _05765_ _05920_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__and3_1
XANTENNA__11029__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13635_ clknet_leaf_77_clk _00748_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ net2346 net232 net431 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
XANTENNA__11631__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12241__A2 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ clknet_leaf_83_clk _00679_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10778_ net1792 net560 net538 _05731_ vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10755__B cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ net1018 _06291_ _06293_ net260 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ clknet_leaf_91_clk _00610_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12448_ cpu.f0.state\[2\] cpu.f0.state\[3\] cpu.f0.state\[7\] net1127 vssd1 vssd1
+ vccd1 vccd1 _06248_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10004__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12379_ net1119 net1850 net529 net1069 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14118_ clknet_leaf_4_clk _01231_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08879__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06940_ net954 cpu.RF0.registers\[11\]\[26\] net775 vssd1 vssd1 vccd1 vccd1 _02231_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_43_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14049_ clknet_leaf_66_clk _01162_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_06871_ net1049 net797 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__and2_1
XANTENNA__11806__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ net304 _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
X_09590_ net494 _04865_ _04879_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__a21o_1
XANTENNA__13805__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ cpu.RF0.registers\[0\]\[6\] net663 net550 vssd1 vssd1 vccd1 vccd1 _03832_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12210__B _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ _03751_ _03754_ _03758_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10011__A cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ cpu.RF0.registers\[29\]\[0\] net601 _02711_ _02712_ _02713_ vssd1 vssd1 vccd1
+ vccd1 _02714_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08119__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13955__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11541__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ net523 _02644_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__nand2_2
XANTENNA__12232__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07958__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08416__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__Q a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06862__C net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07285_ cpu.RF0.registers\[15\]\[7\] net590 _02546_ _02553_ net622 vssd1 vssd1 vccd1
+ vccd1 _02576_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout314_A _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ cpu.RF0.registers\[9\]\[31\] net699 net638 cpu.RF0.registers\[26\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1056_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10952__Y _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 cpu.RF0.registers\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 a1.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10546__A2 a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold242 cpu.RF0.registers\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 cpu.RF0.registers\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold264 cpu.RF0.registers\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13878__RESET_B net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13335__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 _00338_ vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 a1.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout683_A _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 cpu.RF0.registers\[14\]\[8\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _02009_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_8
Xfanout722 _02002_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
X_09926_ net127 _05211_ _05208_ net631 vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout733 cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_4
Xfanout744 _05985_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_2
Xfanout755 _05638_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 net768 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_2
X_09857_ _02004_ _05146_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout850_A _02041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 net779 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net801 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_2
XANTENNA__08372__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13485__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08808_ cpu.RF0.registers\[5\]\[19\] net702 _04096_ _04097_ _04098_ vssd1 vssd1 vccd1
+ vccd1 _04099_ sky130_fd_sc_hd__a2111o_1
X_09788_ net296 net294 _04947_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__mux2_1
XANTENNA__06922__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ _03931_ _03933_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11750_ net1647 net185 net344 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__mux2_1
X_10701_ cpu.LCD0.row_1\[107\] net2526 net897 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ net2119 net173 net353 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XANTENNA__11451__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ clknet_leaf_68_clk _00533_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ net2726 net2185 net907 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12223__A2 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07230__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ net58 net919 vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and2_1
X_13351_ clknet_leaf_80_clk _00464_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08045__B _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ net1478 net555 _06194_ net1370 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10494_ net1520 net919 net750 a1.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 _00167_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ clknet_leaf_20_clk cpu.RU0.next_FetchedInstr\[21\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09927__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ _06114_ _06125_ _06127_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12135__X _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ cpu.LCD0.row_2\[90\] _05983_ _06006_ cpu.LCD0.row_1\[34\] vssd1 vssd1 vccd1
+ vccd1 _06063_ sky130_fd_sc_hd__a22o_1
XANTENNA__14260__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net2162 net209 net418 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__mux2_1
X_12095_ cpu.LCD0.nextState\[1\] cpu.LCD0.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05996_
+ sky130_fd_sc_hd__and2b_2
XANTENNA__13828__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11046_ net2808 net214 net428 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11626__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13978__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12997_ clknet_leaf_35_clk _00186_ net1258 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11948_ net1860 net187 net320 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14667_ net1389 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11879_ net2921 net174 net329 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__mux2_1
XANTENNA__11361__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ clknet_leaf_60_clk _00731_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ clknet_leaf_47_clk _01700_ net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[109\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10225__A1 cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ clknet_leaf_103_clk _00662_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ net974 cpu.RF0.registers\[2\]\[18\] net771 vssd1 vssd1 vccd1 vccd1 _02361_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07641__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14603__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__B _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10006__A cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07972_ cpu.RF0.registers\[31\]\[29\] net686 net635 cpu.RF0.registers\[16\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a22o_1
X_09711_ _04921_ _04944_ _04962_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__or4b_1
X_06923_ net1029 cpu.RF0.registers\[17\]\[26\] net805 vssd1 vssd1 vccd1 vccd1 _02214_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11536__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ net439 _03019_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__and2b_1
X_06854_ net1073 net1066 net1068 net1069 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_39_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12929__Q a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ _03801_ _03803_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nor2_1
X_06785_ cpu.RF0.registers\[31\]\[30\] net687 net654 cpu.RF0.registers\[2\]\[30\]
+ _02060_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout264_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09449__A3 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08524_ net1104 cpu.RF0.registers\[16\]\[6\] net841 vssd1 vssd1 vccd1 vccd1 _03815_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09854__B1 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10947__Y _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ cpu.RF0.registers\[22\]\[8\] net669 net655 cpu.RF0.registers\[2\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout431_A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14133__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07406_ net1048 cpu.RF0.registers\[20\]\[0\] net783 vssd1 vssd1 vccd1 vccd1 _02697_
+ sky130_fd_sc_hd__and3_1
X_08386_ net1089 cpu.RF0.registers\[17\]\[10\] net883 vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_80_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ net1061 cpu.RF0.registers\[31\]\[3\] net829 vssd1 vssd1 vccd1 vccd1 _02628_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10963__X _05860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1340_A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ net980 cpu.RF0.registers\[12\]\[7\] net768 vssd1 vssd1 vccd1 vccd1 _02559_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14283__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout898_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ net1076 cpu.RF0.registers\[16\]\[31\] net841 vssd1 vssd1 vccd1 vccd1 _04298_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12508__A3 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10615__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ net1051 cpu.RF0.registers\[22\]\[10\] net801 vssd1 vssd1 vccd1 vccd1 _02490_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11716__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09385__A2 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
Xfanout541 _05494_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
X_09909_ _05173_ _05174_ _05185_ _05171_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a211o_1
XANTENNA__12875__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout552 _02086_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
Xfanout563 _05641_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_2
Xfanout574 _02187_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 _02173_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11446__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ clknet_leaf_22_clk _00109_ net1173 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout596 _02157_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_8
XANTENNA__09424__B _04705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ clknet_leaf_24_clk _00070_ net1210 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ net1722 net241 net336 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ net1428 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08608__X _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14521_ clknet_leaf_50_clk net2147 net1376 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10455__B2 a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net1857 net255 net344 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11181__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14452_ clknet_leaf_24_clk _01562_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_11664_ net1882 net131 net354 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07598__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13500__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13403_ clknet_leaf_12_clk _00516_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10615_ cpu.LCD0.row_1\[21\] cpu.LCD0.row_1\[29\] net901 vssd1 vssd1 vccd1 vccd1
+ _00245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14383_ clknet_leaf_23_clk _01494_ net1178 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_11595_ net1726 net146 net364 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ clknet_leaf_61_clk _00447_ net1346 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10546_ net1135 a1.ADR_I\[17\] net915 _05660_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__a31o_1
XANTENNA__10592__Y _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[4\] net1247 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[4\] sky130_fd_sc_hd__dfrtp_1
X_10477_ net1415 net923 net748 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a21o_1
XANTENNA__13650__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ cpu.LCD0.row_1\[4\] _06015_ _06021_ cpu.LCD0.row_1\[92\] vssd1 vssd1 vccd1
+ vccd1 _06113_ sky130_fd_sc_hd__a22o_1
X_13196_ clknet_leaf_82_clk _00376_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ cpu.LCD0.row_2\[33\] _06004_ _06009_ cpu.LCD0.row_1\[105\] vssd1 vssd1 vccd1
+ vccd1 _06047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06798__X _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14006__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_94_clk_X clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net2779 _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__o21a_1
XANTENNA__11356__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06958__B _02247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ net2152 net925 net273 _05905_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14588__RESET_B net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13030__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14156__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06570_ cpu.RU0.next_dhit net895 _01950_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__or3b_1
XFILLER_0_73_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10446__B2 a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A2 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08240_ cpu.RF0.registers\[13\]\[14\] net657 _03528_ _03530_ net667 vssd1 vssd1 vccd1
+ vccd1 _03531_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_32_clk_X clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07862__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__A1 cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08171_ net1108 cpu.RF0.registers\[23\]\[20\] net846 vssd1 vssd1 vccd1 vccd1 _03462_
+ sky130_fd_sc_hd__and3_1
XANTENNA_48 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__Y _02271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07122_ cpu.RF0.registers\[23\]\[15\] net613 net579 cpu.RF0.registers\[18\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09349__X _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_X clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07053_ cpu.RF0.registers\[10\]\[19\] net569 _02343_ net624 vssd1 vssd1 vccd1 vccd1
+ _02344_ sky130_fd_sc_hd__a211o_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12898__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12371__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__B1 _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__B2 cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ net947 cpu.RF0.registers\[3\]\[29\] net836 vssd1 vssd1 vccd1 vccd1 _03246_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11266__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_X clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ cpu.RF0.registers\[12\]\[27\] net572 _02194_ _02196_ _02140_ vssd1 vssd1
+ vccd1 vccd1 _02197_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07886_ cpu.RF0.registers\[6\]\[29\] _02175_ net577 cpu.RF0.registers\[28\]\[29\]
+ _03176_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__a221o_1
X_09625_ _03146_ net446 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nor2_1
X_06837_ net970 net832 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout646_A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09556_ _03802_ _04039_ _03771_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a21bo_1
X_06768_ net1088 net864 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and2_4
XANTENNA__13523__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__inv_2
XANTENNA__14649__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1496_A cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09487_ _04399_ _04598_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ cpu.LCD0.cnt_500hz\[5\] cpu.LCD0.cnt_500hz\[4\] cpu.LCD0.cnt_500hz\[7\] cpu.LCD0.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__or4_1
XANTENNA__10988__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ cpu.IM0.address_IM\[9\] net551 _03727_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ cpu.RF0.registers\[8\]\[11\] net708 _03641_ _03643_ _03645_ vssd1 vssd1 vccd1
+ vccd1 _03660_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13673__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ net1126 _01805_ net265 vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__or3_1
XANTENNA__09259__X _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ net1831 net203 net388 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__mux2_1
XANTENNA__07605__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__C1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ _05567_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__nand2_1
XANTENNA__13822__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11030__A cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ cpu.f0.i\[13\] _05503_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__nor2_1
X_13050_ clknet_leaf_52_clk _00230_ net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14029__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12001_ net2064 net233 net312 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__mux2_1
XANTENNA__08566__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08030__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ net625 _04551_ net1022 vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__o21a_1
Xfanout1303 net1306 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
Xfanout1314 net1315 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__clkbuf_4
Xfanout1325 net1326 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09435__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07507__X _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1336 net1342 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1347 net1350 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__clkbuf_4
Xfanout1358 net1363 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13053__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06592__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_8
Xfanout1369 net1371 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14179__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout382 _05925_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_6
X_13952_ clknet_leaf_3_clk _01065_ net1160 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout393 _05923_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12903_ clknet_leaf_26_clk _00092_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13883_ clknet_leaf_14_clk _00996_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11904__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12834_ clknet_leaf_15_clk _00053_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09818__B1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08338__X _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12765_ net1545 net496 net281 net1018 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a22o_1
XANTENNA__08097__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ clknet_leaf_47_clk _01606_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11716_ net2650 net192 net346 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12696_ net2247 cpu.LCD0.row_2\[90\] net1001 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14435_ clknet_leaf_16_clk _01546_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ net1972 net194 net357 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__mux2_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__A1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 gpio_in[12] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
X_14366_ clknet_leaf_58_clk _01479_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11578_ net1576 net202 net363 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__mux2_1
XANTENNA__08514__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06960__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold808 cpu.LCD0.row_2\[47\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13317_ clknet_leaf_18_clk cpu.RU0.next_FetchedData\[24\] net1192 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[24\] sky130_fd_sc_hd__dfrtp_1
X_10529_ net71 net918 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__and2_1
Xhold819 cpu.RF0.registers\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_70_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14297_ clknet_leaf_14_clk _01410_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13248_ clknet_leaf_43_clk _00428_ net1306 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09048__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13179_ clknet_leaf_34_clk _00359_ net1245 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1508 cpu.RF0.registers\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net2914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07791__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1519 cpu.RF0.registers\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net2925 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06688__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ cpu.RF0.registers\[29\]\[20\] net601 net571 cpu.RF0.registers\[12\]\[20\]
+ _03030_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07671_ net1024 cpu.RF0.registers\[30\]\[16\] net761 vssd1 vssd1 vccd1 vccd1 _02962_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11814__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _03173_ net447 vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand2_1
X_06622_ _01757_ _01984_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__or3_1
XANTENNA__12408__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06553_ cpu.DM0.dhit cpu.f0.state\[3\] cpu.f0.state\[0\] net34 _01939_ vssd1 vssd1
+ vccd1 vccd1 _00021_ sky130_fd_sc_hd__a221o_1
X_09341_ _04412_ _04631_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_89_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13696__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__B _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07296__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06484_ cpu.K0.keyvalid _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__nand2_1
X_09272_ net296 _04558_ _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o211a_1
XANTENNA__07835__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08127__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08223_ cpu.RF0.registers\[29\]\[14\] net673 net641 cpu.RF0.registers\[19\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07031__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10954__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_A _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ cpu.RF0.registers\[11\]\[20\] net689 net679 cpu.RF0.registers\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12592__A1 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__Q a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07105_ cpu.RF0.registers\[20\]\[14\] net594 net571 cpu.RF0.registers\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08085_ net1080 cpu.RF0.registers\[20\]\[22\] net874 vssd1 vssd1 vccd1 vccd1 _03376_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_77_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08143__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1136_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ net965 cpu.RF0.registers\[3\]\[19\] net821 vssd1 vssd1 vccd1 vccd1 _02327_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13076__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1303_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14321__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _04275_ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1411_A cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _03218_ _03219_ _03220_ _03221_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14471__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ cpu.RF0.registers\[25\]\[28\] net568 net566 cpu.RF0.registers\[11\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12913__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _04026_ _04471_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10880_ net735 _05140_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ net493 _04775_ _04814_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_17_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08079__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12550_ cpu.f0.state\[5\] _06308_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12280__B1 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ net1504 net236 net372 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _05487_ net257 cpu.f0.i\[10\] vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__a21o_1
XANTENNA__10830__B2 _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14220_ clknet_leaf_79_clk _01333_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11432_ net2335 net136 net382 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08787__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ clknet_leaf_81_clk _01264_ net1291 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10594__A0 cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ net2708 net148 net393 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08251__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13102_ clknet_leaf_53_clk _00282_ net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10314_ net2881 net724 _05554_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__o21a_1
X_14082_ clknet_leaf_94_clk _01195_ net1222 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ net2694 net178 net400 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09736__C1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ clknet_leaf_32_clk _00011_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.DM0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_56_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ net526 net541 _05495_ net725 vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1100 net1108 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1111 cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09751__A2 _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
XANTENNA__13569__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _05438_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__xnor2_1
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_2
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
Xfanout1155 net1167 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1177 net1179 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_4
Xfanout1188 net1190 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_4
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1199 net1211 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_2
X_13935_ clknet_leaf_87_clk _01048_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06795__Y _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08711__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11634__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload5_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_102_clk _00979_ net1215 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10758__B _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07413__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12817_ clknet_leaf_32_clk _00036_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_13797_ clknet_leaf_3_clk _00910_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12748_ cpu.f0.write_data\[6\] net497 _01762_ _01772_ vssd1 vssd1 vccd1 vccd1 _01727_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12271__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07817__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__A1 cpu.IM0.address_IM\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ net2544 net2471 net1007 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08490__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418_ clknet_leaf_31_clk net1616 net1205 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08244__A _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13099__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ clknet_leaf_28_clk _01462_ net1183 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10585__A0 _05680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 cpu.RF0.registers\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14344__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 cpu.RF0.registers\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 a1.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 cpu.FetchedInstr\[15\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 cpu.RF0.registers\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _04198_ _04199_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__or2_1
XANTENNA__11809__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ cpu.IM0.address_IM\[3\] cpu.IM0.address_IM\[2\] cpu.IM0.address_IM\[4\] vssd1
+ vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10713__S net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07147__X _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07202__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ cpu.RF0.registers\[5\]\[16\] net702 _04129_ _04130_ _04131_ vssd1 vssd1 vccd1
+ vccd1 _04132_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10888__A1 _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14494__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1305 cpu.RF0.registers\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07753__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1316 cpu.RF0.registers\[12\]\[5\] vssd1 vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08410__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12936__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1327 cpu.RF0.registers\[25\]\[14\] vssd1 vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ net1095 cpu.RF0.registers\[23\]\[18\] net845 vssd1 vssd1 vccd1 vccd1 _04063_
+ sky130_fd_sc_hd__and3_1
Xhold1338 cpu.RF0.registers\[28\]\[22\] vssd1 vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 a1.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
X_07723_ _03010_ _03011_ _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_85_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__A cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07026__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11544__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _02832_ _02868_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06865__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12937__Q a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06605_ cpu.LCD0.nextState\[2\] net556 _01975_ net1350 vssd1 vssd1 vccd1 vccd1 _01755_
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_88_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07585_ net965 cpu.RF0.registers\[1\]\[12\] net805 vssd1 vssd1 vccd1 vccd1 _02876_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1086_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ net305 _04607_ _04614_ _04480_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06536_ _01895_ _01896_ _01900_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07610__X _02901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10812__A1 cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09255_ net301 _04528_ _04529_ _04385_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__o22a_1
X_06467_ net1130 cpu.RU0.state\[4\] net1409 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout511_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout609_A _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08206_ cpu.RF0.registers\[15\]\[21\] net682 net651 cpu.RF0.registers\[7\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09186_ _04470_ _04476_ net474 vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__mux2_1
X_06398_ net2803 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__inv_2
XANTENNA__07696__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12565__A1 cpu.SR1.char_in\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ cpu.RF0.registers\[13\]\[23\] net659 net638 cpu.RF0.registers\[26\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__a22o_1
XANTENNA__08233__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08068_ _03356_ _03357_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout880_A _02008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07019_ net1066 net633 net519 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1306_X net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07057__X _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ cpu.IM0.address_IM\[15\] _05284_ cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1
+ vccd1 _05307_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ net2037 net186 net316 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__mux2_1
XANTENNA__09497__B2 _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ clknet_leaf_6_clk _00833_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ cpu.DM0.readdata\[30\] _04517_ net734 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__mux2_1
XANTENNA__10500__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14217__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ clknet_leaf_67_clk _00764_ net1298 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ net723 _05244_ _05791_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12602_ cpu.LCD0.row_2\[4\] cpu.SR1.char_in\[4\] net1012 vssd1 vssd1 vccd1 vccd1
+ _01595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13582_ clknet_leaf_1_clk _00695_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10794_ cpu.f0.data_adr\[23\] _04577_ net989 vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ cpu.f0.i\[29\] _06301_ _06303_ net260 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__o211a_1
XANTENNA__10803__B2 _05749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13241__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14367__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ cpu.f0.i\[3\] cpu.f0.i\[4\] _06256_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__and3_1
XANTENNA__12809__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14203_ clknet_leaf_12_clk _01316_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ net1983 net197 net382 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12395_ net1629 cpu.DM0.data_i\[5\] net733 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__mux2_1
XANTENNA__08224__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08999__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14134_ clknet_leaf_71_clk _01247_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ net1871 net212 net392 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
XANTENNA__13391__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06786__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12959__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ clknet_leaf_77_clk _01178_ net1335 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11277_ net2480 net226 net401 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__mux2_1
X_13016_ clknet_leaf_36_clk _00205_ net1260 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
X_10228_ net2870 net726 _05479_ _05481_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 cpu.LCD0.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net630 _04639_ net932 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09623__A _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07499__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ clknet_leaf_84_clk _01031_ net1270 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13849_ clknet_leaf_42_clk _00962_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12244__B1 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ net1054 cpu.RF0.registers\[27\]\[2\] net777 vssd1 vssd1 vccd1 vccd1 _02661_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06982__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08463__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09040_ net1027 cpu.RF0.registers\[21\]\[31\] net795 vssd1 vssd1 vccd1 vccd1 _04331_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09412__A1 _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 cpu.RF0.registers\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09412__B2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold413 cpu.LCD0.row_1\[83\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold424 cpu.RF0.registers\[23\]\[5\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__A2 _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold435 cpu.RF0.registers\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload31_A clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 cpu.RF0.registers\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06777__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold457 cpu.RF0.registers\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 cpu.RF0.registers\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11539__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09942_ _05224_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__or2_1
XANTENNA__12807__RESET_B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold479 cpu.FetchedInstr\[27\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_2
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout915 _01860_ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
Xfanout926 net928 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ cpu.IM0.address_IM\[3\] _02606_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_5_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 net942 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_2
Xfanout948 net950 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 net960 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__buf_2
Xhold1102 cpu.LCD0.row_1\[89\] vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ cpu.RF0.registers\[27\]\[19\] net711 net699 cpu.RF0.registers\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 cpu.RF0.registers\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 cpu.RF0.registers\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 cpu.RF0.registers\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1146 cpu.RF0.registers\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _04045_ _03669_ _03668_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand3b_1
Xhold1157 cpu.RF0.registers\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 cpu.K0.code\[5\] vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06876__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1179 cpu.LCD0.row_2\[58\] vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ net956 cpu.RF0.registers\[9\]\[17\] net756 vssd1 vssd1 vccd1 vccd1 _02997_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08686_ cpu.RF0.registers\[29\]\[1\] net673 _02059_ cpu.RF0.registers\[25\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a22o_1
X_07637_ cpu.RF0.registers\[9\]\[13\] net573 _02920_ _02921_ _02925_ vssd1 vssd1 vccd1
+ vccd1 _02928_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13264__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ cpu.RF0.registers\[27\]\[8\] net591 _02846_ _02849_ _02850_ vssd1 vssd1 vccd1
+ vccd1 _02859_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_76_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ _04595_ _04597_ _04481_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a21bo_1
X_06519_ cpu.f0.num\[22\] net1019 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__or2_1
XANTENNA__10797__A0 cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ cpu.RF0.registers\[4\]\[5\] net587 net575 cpu.RF0.registers\[14\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a22o_1
XANTENNA__08454__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _04369_ _04386_ net454 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11797__X _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ net468 _03729_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_1
XANTENNA__08206__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ net2060 net138 net410 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
X_12180_ cpu.LCD0.row_1\[106\] _06009_ _06011_ cpu.LCD0.row_2\[50\] _06078_ vssd1
+ vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10861__B _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ net1941 net147 net420 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
XANTENNA__10206__X _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 cpu.RF0.registers\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 cpu.RF0.registers\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07228__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ net2072 net158 net426 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08050__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10721__A0 cpu.f0.data_adr\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11184__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13607__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ cpu.RF0.registers\[29\]\[1\] net254 net317 vssd1 vssd1 vccd1 vccd1 _01369_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13703_ clknet_leaf_80_clk _00816_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ net739 _04663_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__nand2_1
X_14683_ net1405 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09890__A1 cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11895_ net2703 net129 net326 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ clknet_leaf_94_clk _00747_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10846_ net723 _05191_ _05779_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13757__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13565_ clknet_leaf_66_clk _00678_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ cpu.IM0.address_IM\[18\] net1014 net285 _05730_ vssd1 vssd1 vccd1 vccd1 _05731_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08445__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10788__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ net1018 _06291_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13496_ clknet_leaf_6_clk _00609_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12447_ net2038 net730 net500 _06247_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__o22a_1
XANTENNA__10004__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08522__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ net1119 net2577 net529 net1072 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11359__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ clknet_leaf_10_clk _01230_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11329_ net2138 net155 net394 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13137__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ clknet_leaf_4_clk _01161_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ net1038 cpu.RF0.registers\[20\]\[27\] net781 vssd1 vssd1 vccd1 vccd1 _02161_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07425__X _02716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07144__Y _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _03821_ _03825_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__or3_2
XANTENNA__14532__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__C _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ cpu.RF0.registers\[12\]\[8\] net697 _03759_ _03760_ _03761_ vssd1 vssd1 vccd1
+ vccd1 _03762_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09881__A1 cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ net972 cpu.RF0.registers\[8\]\[0\] net813 vssd1 vssd1 vccd1 vccd1 _02713_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12217__B1 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12768__B2 cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload79_A clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07353_ cpu.IG0.Instr\[9\] net742 _02208_ net1068 vssd1 vssd1 vccd1 vccd1 _02644_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06862__D net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07284_ _02571_ _02572_ _02573_ _02574_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__nor4_1
XFILLER_0_66_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ cpu.RF0.registers\[15\]\[31\] net682 net646 cpu.RF0.registers\[21\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_57_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout307_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 _01529_ vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold221 cpu.RF0.registers\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 cpu.RF0.registers\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10546__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 cpu.RF0.registers\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 cpu.LCD0.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 cpu.RF0.registers\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold276 cpu.RF0.registers\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 cpu.RF0.registers\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout701 _02022_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_8
X_09925_ _05209_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nor2_1
XANTENNA__09815__X _05106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout712 _02009_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
Xhold298 cpu.RF0.registers\[18\]\[19\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout723 _02001_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
XANTENNA__14062__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_2
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _05980_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_2
Xfanout756 net758 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
X_09856_ _04452_ _05144_ _05145_ _04451_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__o211ai_1
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_2
Xfanout789 _02153_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08807_ net1083 cpu.RF0.registers\[29\]\[19\] net849 vssd1 vssd1 vccd1 vccd1 _04098_
+ sky130_fd_sc_hd__and3_1
X_09787_ _03540_ _05076_ net511 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06999_ net1034 cpu.RF0.registers\[21\]\[23\] net795 vssd1 vssd1 vccd1 vccd1 _02290_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11259__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _04027_ _04028_ _03967_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08669_ cpu.RF0.registers\[10\]\[2\] net692 net686 cpu.RF0.registers\[31\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a22o_1
XANTENNA__11732__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ net2235 cpu.LCD0.row_1\[114\] net897 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07883__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net1936 net193 net353 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10631_ cpu.LCD0.row_1\[37\] cpu.LCD0.row_1\[45\] net900 vssd1 vssd1 vccd1 vccd1
+ _00261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11033__A _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ clknet_leaf_8_clk _00463_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10562_ net1133 net1692 net913 _05668_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ _06075_ _06186_ _06193_ net556 vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13281_ clknet_leaf_20_clk cpu.RU0.next_FetchedInstr\[20\] net1169 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[20\] sky130_fd_sc_hd__dfrtp_1
X_10493_ net1487 net921 net749 a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 _00166_
+ sky130_fd_sc_hd__a22o_1
X_12232_ cpu.LCD0.row_2\[36\] _06004_ _06030_ cpu.LCD0.row_1\[44\] _06128_ vssd1 vssd1
+ vccd1 vccd1 _06129_ sky130_fd_sc_hd__a221o_1
XANTENNA__09927__A2 _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08342__A _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14405__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11179__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net1427 _01965_ _06062_ net1378 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__o211a_1
XANTENNA__09725__X _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ net1865 net202 net419 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
X_12094_ cpu.LCD0.nextState\[5\] cpu.LCD0.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05995_
+ sky130_fd_sc_hd__and2_2
XANTENNA__12799__A cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11907__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11045_ net1995 net217 net426 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__mux2_1
XANTENNA__10811__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14555__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09560__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__A1 cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06913__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__A cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ clknet_leaf_29_clk _00185_ net1202 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__A0 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__A cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ net2361 net189 net318 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__mux2_1
XANTENNA__07124__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11642__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ net1388 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_15_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07874__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11670__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ net2572 net193 net329 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__mux2_1
X_13617_ clknet_leaf_76_clk _00730_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ cpu.DM0.readdata\[0\] net738 net722 vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__o21ai_1
X_14597_ clknet_leaf_49_clk _01699_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[108\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ clknet_leaf_80_clk _00661_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ clknet_leaf_82_clk _00592_ net1284 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14305__RESET_B net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10387__A1_N net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14085__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11089__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__C _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ cpu.RF0.registers\[1\]\[29\] _02007_ net657 cpu.RF0.registers\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09710_ _04899_ _04971_ _04977_ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__and4_1
XANTENNA__11817__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06922_ net543 _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__o21ai_4
XANTENNA__12150__A2 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _04928_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__and2_1
X_06853_ net1049 net806 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13922__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09572_ net494 _04040_ _04847_ _04861_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a311o_2
X_06784_ _02071_ _02072_ _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__or4_1
XANTENNA__10022__A cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08523_ net1103 cpu.RF0.registers\[23\]\[6\] net846 vssd1 vssd1 vccd1 vccd1 _03814_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07034__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07865__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ cpu.RF0.registers\[5\]\[8\] net703 net675 cpu.RF0.registers\[6\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a22o_1
XANTENNA__10464__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07405_ net1048 cpu.RF0.registers\[19\]\[0\] net823 vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07331__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08385_ net1093 cpu.RF0.registers\[26\]\[10\] net860 vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1166_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ net975 cpu.RF0.registers\[4\]\[3\] net782 vssd1 vssd1 vccd1 vccd1 _02627_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13302__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ net1062 cpu.RF0.registers\[18\]\[7\] net772 vssd1 vssd1 vccd1 vccd1 _02558_
+ sky130_fd_sc_hd__and3_1
X_09006_ net934 cpu.RF0.registers\[4\]\[31\] net874 vssd1 vssd1 vccd1 vccd1 _04297_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ net1051 cpu.RF0.registers\[18\]\[10\] net771 vssd1 vssd1 vccd1 vccd1 _02489_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout793_A _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14578__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net521 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_2
Xfanout531 _06221_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ cpu.IM0.address_IM\[6\] _02797_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__xor2_1
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 _05640_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_6
XANTENNA__07506__A cpu.IG0.Instr\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 _02171_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_6
X_09839_ _02604_ _05064_ _04480_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__o21ai_2
Xfanout597 _02155_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_6
XANTENNA__08896__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14400__Q cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ clknet_leaf_31_clk _00069_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11801_ net2514 net247 net336 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ net2539 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11462__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14520_ clknet_leaf_49_clk net2466 net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11732_ net2325 net238 net343 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07241__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14451_ clknet_leaf_24_clk _01561_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_11663_ net2794 net138 net354 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07871__A3 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ clknet_leaf_93_clk _00515_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10614_ cpu.LCD0.row_1\[20\] cpu.LCD0.row_1\[28\] net899 vssd1 vssd1 vccd1 vccd1
+ _00244_ sky130_fd_sc_hd__mux2_1
XANTENNA__12601__A0 cpu.LCD0.row_2\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ clknet_leaf_22_clk _01493_ net1178 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11594_ net2041 net149 net363 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13333_ clknet_leaf_61_clk _00446_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10545_ net48 net916 vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[3\] net1245 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[3\] sky130_fd_sc_hd__dfrtp_1
X_10476_ a1.curr_state\[1\] net1135 a1.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _05642_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_62_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12215_ net1433 net555 _06112_ net1359 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__o211a_1
X_13195_ clknet_leaf_30_clk _00375_ net1208 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ cpu.LCD0.row_2\[9\] _05998_ _06033_ cpu.LCD0.row_2\[73\] _06045_ vssd1 vssd1
+ vccd1 vccd1 _06046_ sky130_fd_sc_hd__a221o_1
XANTENNA__09781__B1 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11637__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ cpu.LCD0.cnt_500hz\[14\] _05978_ _05958_ vssd1 vssd1 vccd1 vccd1 _05979_
+ sky130_fd_sc_hd__a21boi_1
XANTENNA__07139__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ cpu.f0.write_data\[31\] _05904_ net985 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__mux2_1
XANTENNA__08887__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12979_ clknet_leaf_22_clk net1497 net1171 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09836__B2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07847__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08247__A _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07311__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ clknet_leaf_31_clk _01750_ net1206 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_16 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12199__A2 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08170_ net949 cpu.RF0.registers\[1\]\[20\] net885 vssd1 vssd1 vccd1 vccd1 _03461_
+ sky130_fd_sc_hd__and3_1
XANTENNA_38 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09064__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07121_ cpu.RF0.registers\[17\]\[15\] net605 net591 cpu.RF0.registers\[27\]\[15\]
+ _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06822__A1 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07052_ cpu.RF0.registers\[23\]\[19\] net614 net603 cpu.RF0.registers\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XANTENNA__10242__C_N net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__08413__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__09221__C1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07378__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__A1 cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07029__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11547__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09525__B _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ net947 cpu.RF0.registers\[6\]\[29\] net852 vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__and3_1
X_06905_ net1038 cpu.RF0.registers\[30\]\[27\] net762 vssd1 vssd1 vccd1 vccd1 _02196_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07326__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ cpu.RF0.registers\[19\]\[29\] net616 net609 cpu.RF0.registers\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__a22o_1
XANTENNA__10134__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_A _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _04619_ _04620_ _04587_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o21ai_1
X_06836_ net969 net832 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__and2_1
XANTENNA__14100__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ _04831_ _04832_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_56_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06767_ net939 net838 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__and2_4
XFILLER_0_56_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout639_A _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__B net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net507 _03796_ cpu.IM0.address_IM\[7\] net553 vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__07838__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ _04042_ _04044_ _04775_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__or3b_1
X_06698_ net1407 net1131 vssd1 vssd1 vccd1 vccd1 cpu.K0.next_keyvalid sky130_fd_sc_hd__nor2_1
XANTENNA__07699__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07302__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14250__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14298__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ cpu.RF0.registers\[0\]\[9\] net661 net547 vssd1 vssd1 vccd1 vccd1 _03728_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1489_A cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13818__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08368_ cpu.RF0.registers\[28\]\[11\] net705 net648 cpu.RF0.registers\[25\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07319_ net982 cpu.RF0.registers\[6\]\[3\] net802 vssd1 vssd1 vccd1 vccd1 _02610_
+ sky130_fd_sc_hd__and3_1
X_08299_ _03571_ _03587_ _03588_ _03589_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1336_X net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ cpu.f0.i\[22\] _05556_ cpu.f0.i\[23\] vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13968__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__B cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ cpu.f0.i\[13\] _05503_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__and2_1
XANTENNA__06899__X _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__A0 _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ cpu.RF0.registers\[30\]\[4\] net243 net312 vssd1 vssd1 vccd1 vccd1 _01404_
+ sky130_fd_sc_hd__mux2_1
X_10192_ net126 _05455_ _05454_ net630 vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B2 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net1306 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__buf_2
XANTENNA__11457__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1315 net1322 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__clkbuf_4
Xfanout1326 net1331 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__buf_2
XANTENNA__12992__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1337 net1339 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout350 _05933_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_8
Xfanout1348 net1350 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 _05931_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_6
Xfanout1359 net1362 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__clkbuf_4
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_8
X_13951_ clknet_leaf_106_clk _01064_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout383 _05925_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_4
Xfanout394 _05922_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12902_ clknet_leaf_26_clk _00091_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13882_ clknet_leaf_97_clk _00995_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13348__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ clknet_leaf_41_clk _00052_ net1267 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[29\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_9_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__A1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12764_ net1452 net496 net281 net1019 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14503_ clknet_leaf_55_clk _01605_ net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11715_ cpu.RF0.registers\[21\]\[16\] net205 net346 vssd1 vssd1 vccd1 vccd1 _01128_
+ sky130_fd_sc_hd__mux2_1
X_12695_ net2394 net2208 net1009 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XANTENNA__07402__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13498__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ net1658 net198 net354 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__mux2_1
X_14434_ clknet_leaf_16_clk _01545_ net1195 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__A1 _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08254__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14365_ clknet_leaf_57_clk _01478_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput36 gpio_in[13] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_103_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11577_ net1626 net215 net363 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__mux2_1
Xwire773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_2
X_13316_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[23\] net1169 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[23\] sky130_fd_sc_hd__dfrtp_1
X_10528_ net1132 net1604 net913 _05651_ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_2
Xhold809 cpu.RF0.registers\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ clknet_leaf_18_clk _01409_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ clknet_leaf_34_clk _00427_ net1250 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08006__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net8 net752 net562 a1.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13178_ clknet_leaf_34_clk _00358_ net1247 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10364__A1 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11367__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ net745 _05984_ _05996_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__and3_4
XANTENNA__14123__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1509 cpu.RF0.registers\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net2915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07780__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10116__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07670_ net1024 cpu.RF0.registers\[16\]\[16\] net831 vssd1 vssd1 vccd1 vccd1 _02961_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06985__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07532__A2 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14273__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ _01968_ _01986_ _01988_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__o21ai_1
X_09340_ net473 _04487_ _04623_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__a21oi_2
X_06552_ cpu.DM0.dhit cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nand2_8
XANTENNA__12274__D1 _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ net302 _04401_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06483_ _01867_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08222_ _03407_ _03442_ _03512_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_60_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload61_A clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12865__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08245__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ cpu.RF0.registers\[22\]\[20\] net669 net660 cpu.RF0.registers\[30\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07104_ cpu.RF0.registers\[8\]\[14\] net612 net604 cpu.RF0.registers\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
XANTENNA__07599__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12592__A2 _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08084_ _03339_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07035_ net963 cpu.RF0.registers\[7\]\[19\] net816 vssd1 vssd1 vccd1 vccd1 _02326_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1031_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08440__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _02250_ _03148_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07937_ cpu.RF0.registers\[24\]\[30\] net608 _03227_ net621 vssd1 vssd1 vccd1 vccd1
+ _03228_ sky130_fd_sc_hd__a211o_1
XANTENNA__14616__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout756_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07868_ _03152_ _03154_ _03156_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or4_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ _04025_ net295 _04402_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a21oi_1
X_06819_ _02108_ _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ net1032 cpu.RF0.registers\[20\]\[22\] net780 vssd1 vssd1 vccd1 vccd1 _03090_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09538_ net277 _04826_ _04828_ _04819_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a211o_1
XANTENNA__13640__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08318__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _03534_ net442 net466 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _05765_ _05766_ net504 vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__and3_1
X_12480_ _05485_ _06268_ _06270_ net263 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_43_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09028__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_clk_X clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08615__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ cpu.RF0.registers\[12\]\[29\] net141 net384 vssd1 vssd1 vccd1 vccd1 _00853_
+ sky130_fd_sc_hd__mux2_1
X_14150_ clknet_leaf_5_clk _01263_ net1145 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ net1874 net156 net390 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ clknet_leaf_51_clk net2706 net1379 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08053__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ net527 _05551_ _05552_ _05553_ net728 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a311o_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ clknet_leaf_63_clk _01194_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14146__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ net2269 _05827_ net398 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13032_ clknet_leaf_55_clk _00004_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10244_ cpu.f0.i\[10\] _05487_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07747__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1101 net1108 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
Xfanout1112 cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10175_ _05419_ _05439_ _05429_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__o21a_1
Xfanout1123 cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_2
Xfanout1134 _01790_ vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_31_clk_X clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1145 net1148 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_4
Xfanout1156 net1167 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14296__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1167 net1211 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_2
Xfanout180 _05829_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06970__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
XANTENNA__11915__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13934_ clknet_leaf_0_clk _01047_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__X _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ clknet_leaf_103_clk _00978_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_X clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12816_ clknet_leaf_39_clk _00035_ net1254 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13796_ clknet_leaf_96_clk _00909_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08475__B1 cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ cpu.f0.i\[6\] _01871_ _06345_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11650__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12678_ net2724 net2352 net1009 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XANTENNA__10821__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14417_ clknet_leaf_32_clk _01528_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11629_ net1691 net141 net360 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_104_clk_X clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09975__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ clknet_leaf_27_clk _01461_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10585__A1 cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold606 cpu.RF0.registers\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold617 cpu.RF0.registers\[18\]\[8\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 cpu.RF0.registers\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ clknet_leaf_81_clk _01392_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold639 cpu.RF0.registers\[27\]\[22\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10337__A1 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14639__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11097__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08840_ net1075 cpu.RF0.registers\[28\]\[16\] net867 vssd1 vssd1 vccd1 vccd1 _04131_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07753__A2 _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1306 cpu.DM0.readdata\[8\] vssd1 vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1317 cpu.RF0.registers\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ net948 cpu.RF0.registers\[13\]\[18\] net850 vssd1 vssd1 vccd1 vccd1 _04062_
+ sky130_fd_sc_hd__and3_1
Xhold1328 cpu.RF0.registers\[23\]\[4\] vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06961__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1339 cpu.RF0.registers\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11825__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ cpu.RF0.registers\[16\]\[17\] net582 _02990_ _02997_ _03004_ vssd1 vssd1
+ vccd1 vccd1 _03013_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13663__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09091__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _02410_ _02436_ _02903_ _02940_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_81_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06604_ cpu.LCD0.currentState\[2\] net555 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_66_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07584_ net1046 cpu.RF0.registers\[20\]\[12\] net781 vssd1 vssd1 vccd1 vccd1 _02875_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14019__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09323_ _04485_ _04606_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__nor2_1
X_06535_ _01897_ _01903_ _01907_ _01918_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__or4_1
XANTENNA__07042__C net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11560__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_A _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _04482_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1079_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ _01861_ _01863_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__nand2_1
XANTENNA__10812__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08205_ cpu.RF0.registers\[29\]\[21\] net672 _03483_ _03486_ _03488_ vssd1 vssd1
+ vccd1 vccd1 _03496_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06881__C net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__Q a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09185_ _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06397_ net1019 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14169__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1246_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ cpu.RF0.registers\[5\]\[23\] net702 net636 cpu.RF0.registers\[16\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10576__A1 cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12391__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ cpu.RF0.registers\[9\]\[25\] net701 net648 cpu.RF0.registers\[25\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__a22o_1
XANTENNA__10904__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13193__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ cpu.RF0.registers\[0\]\[23\] net617 _02304_ _02308_ vssd1 vssd1 vccd1 vccd1
+ _02309_ sky130_fd_sc_hd__o22a_2
XANTENNA__08170__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07744__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ cpu.RF0.registers\[22\]\[26\] net670 net638 cpu.RF0.registers\[26\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11735__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ net1869 net189 net314 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__mux2_1
XANTENNA__12420__A cpu.DM0.data_i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net2764 net142 net431 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__mux2_1
XANTENNA__07514__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10500__B2 a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ cpu.DM0.readdata\[10\] net738 net722 vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__o21a_1
X_13650_ clknet_leaf_61_clk _00763_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12601_ cpu.LCD0.row_2\[3\] net1552 net1012 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__mux2_1
X_13581_ clknet_leaf_101_clk _00694_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ net2936 net558 net536 _05742_ vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11470__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12532_ cpu.f0.i\[29\] _06301_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10803__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12863__Q cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ _06258_ _06259_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14202_ clknet_leaf_93_clk _01315_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11414_ net1945 net208 net382 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12394_ net2798 cpu.DM0.data_i\[4\] net733 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_73_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13536__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ clknet_leaf_73_clk _01246_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11345_ net1948 net219 net390 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
XANTENNA__10814__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14064_ clknet_leaf_75_clk _01177_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ net2406 net230 net401 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13015_ clknet_leaf_43_clk _00204_ net1303 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
X_10227_ net528 net309 net1021 vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ net126 _05424_ _05421_ net630 vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a211o_1
Xhold3 cpu.RU0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11645__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11819__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ cpu.IM0.address_IM\[21\] _03078_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__B net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13917_ clknet_leaf_88_clk _01030_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08696__B1 _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_7_clk _00961_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08448__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__B2 cpu.LCD0.row_2\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__B1_N net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ clknet_leaf_68_clk _00892_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11380__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14311__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07120__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07797__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__B1 cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10558__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08542__X _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09412__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14461__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 cpu.RF0.registers\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _00307_ vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10724__S net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 cpu.RF0.registers\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold436 cpu.RF0.registers\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12903__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold447 cpu.FetchedInstr\[26\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold458 cpu.RF0.registers\[15\]\[17\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ cpu.IG0.Instr\[29\] cpu.IM0.address_IM\[9\] net520 vssd1 vssd1 vccd1 vccd1
+ _05225_ sky130_fd_sc_hd__and3_1
Xhold469 cpu.RF0.registers\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06503__A cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload24_A clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout905 _01940_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08421__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_5_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ cpu.IM0.address_IM\[3\] _02606_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__and2_1
Xfanout938 net942 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_2
XANTENNA__12180__B1 _06011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _00313_ vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ cpu.RF0.registers\[20\]\[19\] net710 net691 cpu.RF0.registers\[10\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07037__C net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1114 cpu.RF0.registers\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 cpu.LCD0.row_2\[38\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11555__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1136 cpu.DM0.readdata\[26\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03699_ _03700_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__xnor2_1
Xhold1147 cpu.RF0.registers\[5\]\[28\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1158 cpu.LCD0.row_1\[82\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 cpu.RF0.registers\[4\]\[1\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ net1033 cpu.RF0.registers\[24\]\[17\] net811 vssd1 vssd1 vccd1 vccd1 _02996_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07334__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12948__Q a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08687__B1 _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ cpu.RF0.registers\[11\]\[1\] net689 net639 cpu.RF0.registers\[26\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_92_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout454_A _02756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10398__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13409__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ net964 cpu.RF0.registers\[14\]\[13\] net764 vssd1 vssd1 vccd1 vccd1 _02927_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08439__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ cpu.RF0.registers\[12\]\[8\] net571 _02837_ _02843_ _02844_ vssd1 vssd1 vccd1
+ vccd1 _02858_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_53_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11290__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _04484_ _04581_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__nand2_1
X_06518_ cpu.f0.num\[7\] net1021 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07498_ _02785_ _02786_ _02787_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__or4_2
XANTENNA__10797__A1 _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13559__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _04373_ _04388_ net449 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
X_06449_ _01826_ _01834_ _01855_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[5\] sky130_fd_sc_hd__and3b_1
XFILLER_0_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ _04457_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout990_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ net935 cpu.RF0.registers\[3\]\[23\] net835 vssd1 vssd1 vccd1 vccd1 _03410_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _04385_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__or2_1
X_11130_ net1916 net149 net419 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
Xhold970 cpu.LCD0.row_2\[9\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 cpu.RF0.registers\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14403__Q cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ net2730 net161 net427 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
Xhold992 cpu.RF0.registers\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12171__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ cpu.IM0.address_IM\[15\] _02434_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__nand2_1
XANTENNA__07717__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10721__A1 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__Q cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11963_ net1758 net237 net316 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10485__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14334__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ clknet_leaf_5_clk _00815_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net2103 net178 net431 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ net1404 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
X_11894_ net2197 net137 net326 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09890__A2 cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10845_ cpu.DM0.readdata\[5\] net738 net722 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__o21a_1
XANTENNA__11029__A2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13633_ clknet_leaf_63_clk _00746_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10776_ cpu.f0.data_adr\[18\] _05117_ net991 vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__mux2_1
X_13564_ clknet_leaf_8_clk _00677_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10788__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__B2 cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14484__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12515_ _06291_ _06292_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__nor2_1
XANTENNA__07410__C net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ clknet_leaf_64_clk _00608_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10892__X _05814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12926__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12446_ cpu.DM0.data_i\[31\] net534 vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08803__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ net1120 net1468 net530 net1079 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ net2750 net160 net395 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
X_14116_ clknet_leaf_95_clk _01229_ net1219 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14047_ clknet_leaf_0_clk _01160_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11259_ net2589 net154 net402 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11375__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__B _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12465__A1 cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08669__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12210__D _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08470_ net946 cpu.RF0.registers\[9\]\[8\] net863 vssd1 vssd1 vccd1 vccd1 _03761_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09881__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ net972 cpu.RF0.registers\[3\]\[0\] net823 vssd1 vssd1 vccd1 vccd1 _02712_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13701__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10228__B1 _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07352_ net524 _02641_ _02607_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12768__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08416__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07283_ cpu.RF0.registers\[14\]\[7\] net575 _02556_ _02558_ _02563_ vssd1 vssd1 vccd1
+ vccd1 _02574_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09022_ _04309_ _04310_ _04311_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09809__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold200 cpu.RF0.registers\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 a1.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__Y _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 cpu.RF0.registers\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 cpu.SR1.char_in\[1\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 cpu.RF0.registers\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 cpu.RF0.registers\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14207__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold266 cpu.RF0.registers\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 a1.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 cpu.FetchedInstr\[22\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ cpu.IM0.address_IM\[6\] _05189_ cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1
+ vccd1 _05210_ sky130_fd_sc_hd__a21oi_1
Xhold299 cpu.c0.count\[13\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net704 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_6
Xfanout713 _02007_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_8
Xfanout724 net726 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1111_A cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12153__B1 _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_2
Xfanout746 _05980_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _04452_ _05144_ _05145_ _04451_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__o211a_4
XANTENNA__07990__C net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net758 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__buf_4
XANTENNA_fanout571_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _02181_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11285__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 _02164_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout669_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__A3 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net1086 cpu.RF0.registers\[19\]\[19\] net836 vssd1 vssd1 vccd1 vccd1 _04097_
+ sky130_fd_sc_hd__and3_1
X_09786_ _03540_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__nor2_1
X_06998_ net1035 cpu.RF0.registers\[22\]\[23\] net799 vssd1 vssd1 vccd1 vccd1 _02289_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07064__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12456__A1 cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ _03964_ _03966_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_65_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_X net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ cpu.RF0.registers\[1\]\[2\] net713 net675 cpu.RF0.registers\[6\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a22o_1
XANTENNA__13887__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__X _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ net1045 cpu.RF0.registers\[29\]\[13\] net792 vssd1 vssd1 vccd1 vccd1 _02910_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ cpu.RF0.registers\[5\]\[4\] net703 net655 cpu.RF0.registers\[2\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12949__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ cpu.LCD0.row_1\[36\] cpu.LCD0.row_1\[44\] net903 vssd1 vssd1 vccd1 vccd1
+ _00260_ sky130_fd_sc_hd__mux2_1
XANTENNA__12759__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ net57 net920 vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08293__D1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07230__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _05982_ net744 _05996_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13280_ clknet_leaf_21_clk cpu.RU0.next_FetchedInstr\[19\] net1176 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[19\] sky130_fd_sc_hd__dfrtp_1
X_10492_ net1502 net916 net751 a1.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 _00165_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08623__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ cpu.LCD0.row_1\[12\] _05994_ _06036_ cpu.LCD0.row_1\[20\] vssd1 vssd1 vccd1
+ vccd1 _06128_ sky130_fd_sc_hd__a22o_1
XANTENNA__09388__A1 _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ _06044_ _06046_ _06048_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_9_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07239__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08061__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ net2923 net213 net420 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__mux2_1
X_12093_ net745 _05989_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__and3_4
XANTENNA__12144__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__A _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ net1723 net221 net428 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A1 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09173__B _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10170__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13724__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07405__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ clknet_leaf_35_clk _00184_ net1258 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_56_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11923__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__A1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__B1 _05640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11946_ net2460 net206 net318 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07702__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14665_ cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11877_ net1597 net200 net326 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13874__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ clknet_leaf_75_clk _00729_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10828_ _01852_ _05005_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nor2_1
X_14596_ clknet_leaf_46_clk net2150 net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08823__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ clknet_leaf_92_clk _00660_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10759_ net987 cpu.f0.data_adr\[13\] vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13104__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13478_ clknet_leaf_6_clk _00591_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10274__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ cpu.DM0.readdata\[22\] net730 net500 _06238_ vssd1 vssd1 vccd1 vccd1 _01538_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07929__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__D _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _03257_ _03258_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__or4_1
XANTENNA__13254__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ net525 _02207_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__or2_1
XANTENNA__10146__C1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ _02383_ net441 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__xor2_1
X_06852_ net1069 net1067 net1065 net1072 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__nor4b_2
X_09571_ net277 _04859_ _04852_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a21bo_1
X_06783_ cpu.RF0.registers\[3\]\[30\] net642 net638 cpu.RF0.registers\[26\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_47_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10449__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11833__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ net1104 cpu.RF0.registers\[24\]\[6\] net871 vssd1 vssd1 vccd1 vccd1 _03813_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkload91_A clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ cpu.RF0.registers\[13\]\[8\] net657 _03741_ _03742_ _03743_ vssd1 vssd1 vccd1
+ vccd1 _03744_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07404_ net1048 cpu.RF0.registers\[16\]\[0\] net832 vssd1 vssd1 vccd1 vccd1 _02695_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09067__A0 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ net1090 cpu.RF0.registers\[20\]\[10\] net875 vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_34_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07335_ net1063 cpu.RF0.registers\[19\]\[3\] net824 vssd1 vssd1 vccd1 vccd1 _02626_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12610__A1 cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12664__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1061_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07266_ net1062 cpu.RF0.registers\[31\]\[7\] net829 vssd1 vssd1 vccd1 vccd1 _02557_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08443__A _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09005_ net1076 cpu.RF0.registers\[20\]\[31\] net874 vssd1 vssd1 vccd1 vccd1 _04296_
+ sky130_fd_sc_hd__and3_1
X_07197_ net968 cpu.RF0.registers\[10\]\[10\] net787 vssd1 vssd1 vccd1 vccd1 _02488_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1326_A net1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10924__A1 _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14086__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__B2 _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10912__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 _02209_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09907_ _05193_ _05194_ cpu.IM0.address_IM\[5\] cpu.IM0.pc_enable vssd1 vssd1 vccd1
+ vccd1 _00028_ sky130_fd_sc_hd__o2bb2a_1
Xfanout532 _05848_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_4
Xfanout543 net546 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_6
XANTENNA__13747__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 _02086_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _02195_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_8
Xfanout576 _02184_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_6
X_09838_ _04536_ _04567_ _05124_ _05125_ _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a2111oi_1
Xfanout587 _02171_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_4
Xfanout598 _02155_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_4
X_09769_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__and2b_1
XANTENNA__07225__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ net1698 net251 net337 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__mux2_1
XANTENNA__13897__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12780_ net1572 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07305__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09213__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07522__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ net506 _05912_ _05915_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14450_ clknet_leaf_31_clk _01560_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13127__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11662_ net1870 net140 net356 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08056__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13401_ clknet_leaf_65_clk _00514_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10613_ net2428 net2303 net899 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
X_11593_ net1711 net157 net362 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__mux2_1
X_14381_ clknet_leaf_23_clk _01492_ net1178 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10544_ net1135 a1.ADR_I\[16\] net915 _05659_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13332_ clknet_leaf_61_clk _00445_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08353__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[2\] net1245 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13277__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net26 net752 net562 net2868 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12365__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14522__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ _06102_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__or2_1
X_13194_ clknet_leaf_30_clk _00374_ net1208 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08640__X _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ cpu.LCD0.row_2\[89\] _05983_ _06011_ cpu.LCD0.row_2\[49\] vssd1 vssd1 vccd1
+ vccd1 _06045_ sky130_fd_sc_hd__a22o_1
XANTENNA__09781__A1 _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12076_ _05978_ net502 _05977_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__and3b_1
XFILLER_0_40_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11027_ _04357_ net532 net282 vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10123__A cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11653__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ clknet_leaf_35_clk net1521 net1258 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
X_11929_ net505 _05766_ _05906_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and3_4
XANTENNA__10300__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14648_ clknet_leaf_24_clk _01749_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14052__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ clknet_leaf_54_clk net2375 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07120_ cpu.RF0.registers\[16\]\[15\] net581 net573 cpu.RF0.registers\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08272__A1 cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07051_ _02338_ _02339_ _02340_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_11_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11828__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12513__A cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07783__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07953_ net947 cpu.RF0.registers\[2\]\[29\] net853 vssd1 vssd1 vccd1 vccd1 _03244_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08327__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ net1057 net763 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__and2_4
X_07884_ cpu.RF0.registers\[17\]\[29\] net606 net598 cpu.RF0.registers\[13\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _04360_ _04912_ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__and3_1
X_06835_ net1072 net1069 net1067 net1065 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nor4_1
XANTENNA__11563__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net302 _04844_ _04843_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__o21ba_1
X_06766_ net946 net845 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08505_ cpu.RF0.registers\[0\]\[7\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03796_
+ sky130_fd_sc_hd__o21ai_1
X_09485_ _04041_ _04775_ _04044_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__a21bo_1
X_06697_ net1131 vssd1 vssd1 vccd1 vccd1 cpu.K0.next_state sky130_fd_sc_hd__inv_2
XFILLER_0_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ _03718_ _03719_ _03723_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12394__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ _03654_ _03655_ _03656_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__A0 cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14545__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ net975 cpu.RF0.registers\[8\]\[3\] net813 vssd1 vssd1 vccd1 vccd1 _02609_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09269__A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ cpu.RF0.registers\[20\]\[13\] net710 net642 cpu.RF0.registers\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10070__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ cpu.RF0.registers\[4\]\[9\] net586 _02517_ _02528_ net621 vssd1 vssd1 vccd1
+ vccd1 _02540_ sky130_fd_sc_hd__a2111o_1
X_10260_ _05508_ _05505_ net725 cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1 _00067_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__A1 _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ cpu.IM0.address_IM\[29\] _05443_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__clkbuf_4
Xfanout1316 net1322 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07517__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1327 net1331 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _05936_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_6
Xfanout1338 net1339 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09515__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1349 net1350 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__clkbuf_4
Xfanout351 _05933_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout362 _05930_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_6
X_13950_ clknet_leaf_83_clk _01063_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout373 _05928_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_4
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
Xfanout395 _05922_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12901_ clknet_leaf_26_clk _00090_ net1183 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12569__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13881_ clknet_leaf_14_clk _00994_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11473__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ clknet_leaf_41_clk _00051_ net1267 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[28\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__09279__A0 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14075__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12763_ cpu.f0.write_data\[21\] net498 net279 cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1
+ _01742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14502_ clknet_leaf_45_clk _01604_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[13\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10833__A0 cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11714_ net2782 net176 net348 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12694_ net2513 net2359 net1010 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14433_ clknet_leaf_17_clk _01544_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ net1569 net210 net354 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ clknet_leaf_58_clk _01477_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_5_clk_X clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ net2177 net217 net362 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__mux2_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 gpio_in[14] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08514__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[22\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[22\] sky130_fd_sc_hd__dfrtp_1
X_10527_ net70 net920 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire774 _02172_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_2
X_14295_ clknet_leaf_64_clk _01408_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire785 _02159_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10118__A cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ clknet_leaf_43_clk _00426_ net1304 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ net7 net755 _05640_ a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08811__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11010__A0 cpu.f0.write_data\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13177_ clknet_leaf_34_clk _00357_ net1247 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10389_ _01796_ net270 _05612_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09626__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ cpu.LCD0.row_2\[40\] _06027_ _06028_ cpu.LCD0.row_1\[112\] vssd1 vssd1 vccd1
+ vccd1 _06029_ sky130_fd_sc_hd__a22o_1
X_12059_ net2500 _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10116__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14418__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _01756_ _01977_ _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__or3_1
X_06551_ cpu.f0.state\[5\] _01872_ _01891_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_83_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13442__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14568__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ net434 net288 _04560_ _04559_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a31o_1
X_06482_ _01868_ cpu.K0.code\[3\] cpu.K0.code\[2\] vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__or3b_2
XANTENNA__07296__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08221_ _03477_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10727__S net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ cpu.RF0.registers\[10\]\[20\] net692 net644 cpu.RF0.registers\[3\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__a22o_1
XANTENNA__08245__A1 _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload54_A clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ cpu.RF0.registers\[29\]\[14\] net601 net566 cpu.RF0.registers\[11\]\[14\]
+ _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08083_ _03372_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_9_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07034_ net1040 cpu.RF0.registers\[29\]\[19\] net792 vssd1 vssd1 vccd1 vccd1 _02325_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_77_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11558__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06879__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout484_A _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ cpu.RF0.registers\[5\]\[30\] net603 net573 cpu.RF0.registers\[9\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14098__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ cpu.RF0.registers\[8\]\[28\] net612 net592 cpu.RF0.registers\[27\]\[28\]
+ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a221o_1
XANTENNA__11293__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _04742_ _04807_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13242__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06818_ cpu.CU0.bit30 _02103_ _02107_ _02093_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07798_ net957 cpu.RF0.registers\[4\]\[22\] net781 vssd1 vssd1 vccd1 vccd1 _03089_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07072__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net303 _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__nor2_1
X_06749_ net936 cpu.RF0.registers\[6\]\[30\] net851 vssd1 vssd1 vccd1 vccd1 _02040_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ net300 _04158_ net463 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__mux2_1
XANTENNA__12280__A2 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07800__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08419_ net935 cpu.RF0.registers\[13\]\[9\] net848 vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09399_ net453 _04511_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ net2047 net145 net385 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14406__Q cpu.DM0.readdata\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ net2046 net161 net392 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
XANTENNA__08787__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06798__A1 cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ clknet_leaf_50_clk net2371 net1382 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_10312_ cpu.f0.i\[20\] _05544_ _05550_ net307 vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__o211a_1
XANTENNA__09286__X _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07995__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06798__B2 _02081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14080_ clknet_leaf_2_clk _01193_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11292_ cpu.RF0.registers\[8\]\[22\] net163 net398 vssd1 vssd1 vccd1 vccd1 _00718_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10880__B _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ cpu.f0.i\[10\] _05487_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13031_ clknet_leaf_55_clk _00003_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09736__B2 _04397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10346__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__B1 _06332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1102 net1104 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13315__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ cpu.IM0.address_IM\[27\] _02211_ _02248_ cpu.IM0.address_IM\[26\] vssd1 vssd1
+ vccd1 vccd1 _05439_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1113 cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_1
Xfanout1124 net1127 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_2
Xfanout1135 _01790_ vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_2
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
Xfanout1157 net1158 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_4
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
Xfanout1168 net1170 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_2
Xfanout181 net184 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout192 _05812_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
X_13933_ clknet_leaf_101_clk _01046_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13465__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13864_ clknet_leaf_99_clk _00977_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08078__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ clknet_leaf_39_clk _00034_ net1254 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07413__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13795_ clknet_leaf_79_clk _00908_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11931__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12746_ cpu.f0.write_data\[5\] net497 _01770_ _01771_ vssd1 vssd1 vccd1 vccd1 _01726_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07278__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__B2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08806__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12677_ net2251 net2141 net1002 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ clknet_leaf_32_clk _01527_ net1249 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14118__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11628_ net2369 net144 net361 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__mux2_1
XANTENNA__09975__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ clknet_leaf_28_clk _01460_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11559_ net2651 net159 net367 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold607 cpu.RF0.registers\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 cpu.RF0.registers\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 cpu.f0.num\[14\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09637__A _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14278_ clknet_leaf_5_clk _01391_ net1145 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10790__B _04617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ clknet_leaf_45_clk _00409_ net1312 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07738__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14240__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13753__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1307 cpu.LCD0.row_2\[14\] vssd1 vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 cpu.LCD0.row_2\[80\] vssd1 vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13808__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ cpu.RF0.registers\[10\]\[18\] net693 net644 cpu.RF0.registers\[3\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1329 cpu.RF0.registers\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
X_07721_ cpu.RF0.registers\[14\]\[17\] net576 _02994_ _03003_ _03007_ vssd1 vssd1
+ vccd1 vccd1 _03012_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_85_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12002__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__C net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ _01974_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13958__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07583_ net964 cpu.RF0.registers\[8\]\[12\] net812 vssd1 vssd1 vccd1 vccd1 _02874_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07323__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11841__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06534_ _01919_ _01920_ _01921_ _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__or4_1
X_09322_ _04504_ net272 _04566_ _04463_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07620__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__inv_2
XANTENNA__10273__B2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ net479 _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ cpu.RF0.registers\[5\]\[21\] net704 net671 cpu.RF0.registers\[23\]\[21\]
+ _03494_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09184_ _04471_ _04474_ net458 vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06396_ cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ _03422_ _03423_ _03424_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__nor4_1
XANTENNA__12672__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07977__B1 _03266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ cpu.RF0.registers\[31\]\[25\] net686 _03346_ _03351_ _03355_ vssd1 vssd1
+ vccd1 vccd1 _03357_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13338__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout699_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07017_ _02299_ _02305_ _02306_ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__or4_1
XANTENNA__11288__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07067__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A _02019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13488__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ net936 cpu.RF0.registers\[8\]\[26\] net870 vssd1 vssd1 vccd1 vccd1 _04259_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07919_ net1030 cpu.RF0.registers\[25\]\[30\] net758 vssd1 vssd1 vccd1 vccd1 _03210_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08154__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ cpu.RF0.registers\[2\]\[17\] net654 _04167_ _04171_ _04177_ vssd1 vssd1 vccd1
+ vccd1 _04190_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_19_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ _05455_ _05840_ net721 vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__mux2_4
XFILLER_0_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10500__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10861_ net740 _04830_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nand2_1
XANTENNA__07233__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11751__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ cpu.LCD0.row_2\[2\] cpu.SR1.char_in\[2\] net1000 vssd1 vssd1 vccd1 vccd1
+ _01593_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13580_ clknet_leaf_88_clk _00693_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10792_ net284 _05740_ _05741_ net1013 cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1
+ vccd1 _05742_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_26_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06468__B1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ cpu.f0.i\[28\] _06299_ _06302_ net260 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_26_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14113__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12462_ cpu.f0.i\[3\] _06256_ net261 vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07680__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08064__C net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201_ clknet_leaf_42_clk _01314_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11413_ net1890 net203 net385 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13040__Q cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12582__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ net1710 cpu.DM0.data_i\[3\] net733 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14132_ clknet_leaf_71_clk _01245_ net1339 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11344_ net1845 net221 net392 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14263__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11198__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09176__B _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14063_ clknet_leaf_83_clk _01176_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ net1940 net233 net400 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ clknet_leaf_43_clk _00203_ net1303 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
X_10226_ cpu.f0.data_adr\[8\] net725 _05480_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08393__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10157_ _05422_ _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 _00016_ vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07705__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ cpu.IM0.address_IM\[21\] _03078_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08145__B1 cpu.IM0.address_IM\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__C1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13916_ clknet_leaf_12_clk _01029_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07499__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13847_ clknet_leaf_66_clk _00960_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11661__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12244__A2 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ clknet_leaf_60_clk _00891_ net1344 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__B1 a1.WRITE_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12729_ cpu.f0.state\[7\] cpu.f0.state\[5\] _06317_ vssd1 vssd1 vccd1 vccd1 _01760_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14606__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A1 _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08605__D1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10558__A2 a1.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11755__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold404 cpu.RF0.registers\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13934__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 cpu.RF0.registers\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 cpu.RF0.registers\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 cpu.RF0.registers\[21\]\[19\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 cpu.RF0.registers\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ cpu.IG0.Instr\[29\] net520 cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1
+ _05224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold459 cpu.RF0.registers\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13630__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
Xfanout917 net924 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_2
X_09871_ cpu.IM0.address_IM\[2\] _01787_ _05161_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a21o_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07318__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout939 net941 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_2
XANTENNA_clkload17_A clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _04109_ _04110_ _04111_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_87_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 cpu.RF0.registers\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12521__A cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1115 cpu.RF0.registers\[24\]\[5\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 _01629_ vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 cpu.RF0.registers\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07615__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _03668_ _03669_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_92_clk_X clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1148 cpu.RF0.registers\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13780__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 _00306_ vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07704_ net954 cpu.RF0.registers\[3\]\[17\] net820 vssd1 vssd1 vccd1 vccd1 _02995_
+ sky130_fd_sc_hd__and3_1
X_08684_ cpu.RF0.registers\[3\]\[1\] net644 _03973_ _03974_ vssd1 vssd1 vccd1 vccd1
+ _03975_ sky130_fd_sc_hd__a211o_1
XANTENNA__09830__A _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07635_ net1045 cpu.RF0.registers\[30\]\[13\] net762 vssd1 vssd1 vccd1 vccd1 _02926_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12816__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14136__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout447_A _03300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08439__A1 _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ cpu.RF0.registers\[26\]\[8\] net599 _02840_ _02841_ _02852_ vssd1 vssd1 vccd1
+ vccd1 _02857_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_18_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07988__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ net480 _04593_ _04594_ _04440_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__B2 cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06517_ cpu.f0.num\[5\] _01795_ cpu.f0.num\[3\] _01793_ vssd1 vssd1 vccd1 vccd1 _01906_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ cpu.RF0.registers\[29\]\[5\] net601 _02765_ _02767_ _02780_ vssd1 vssd1 vccd1
+ vccd1 _02788_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1356_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ net478 _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nor2_1
X_06448_ cpu.c0.count\[4\] _01824_ cpu.c0.count\[5\] vssd1 vssd1 vccd1 vccd1 _01855_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13160__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14286__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09939__A1 cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06379_ cpu.f0.num\[6\] vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__inv_2
X_09167_ net468 _03797_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ net1078 cpu.RF0.registers\[18\]\[23\] net855 vssd1 vssd1 vccd1 vccd1 _03409_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _04386_ _04388_ net454 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__C _02019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08049_ _03339_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__inv_2
XANTENNA__10216__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold960 _00265_ vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 cpu.RF0.registers\[26\]\[20\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold982 cpu.RF0.registers\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net1938 net178 net429 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
Xhold993 cpu.LCD0.row_2\[67\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ cpu.IM0.address_IM\[15\] _02434_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__nor2_1
XANTENNA__10182__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_X clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ net505 _05766_ _05910_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_4
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08059__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ clknet_leaf_102_clk _00814_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10913_ _05401_ _05828_ net721 vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__mux2_2
XFILLER_0_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14681_ net1403 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_11893_ net1668 net141 net328 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11481__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ clknet_leaf_4_clk _00745_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10844_ net740 _05073_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nand2_1
XANTENNA__08356__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13503__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07260__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14629__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13563_ clknet_leaf_12_clk _00676_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10775_ a1.ADR_I\[17\] net558 net536 _05729_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09739__X _05030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ _01814_ _06290_ net262 vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__a21bo_1
X_13494_ clknet_leaf_59_clk _00607_ net1348 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12445_ net1750 net731 net501 _06246_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__o22a_1
XANTENNA__13653__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ net1121 net2893 net530 cpu.IG0.Instr\[18\] vssd1 vssd1 vccd1 vccd1 _01502_
+ sky130_fd_sc_hd__a22o_1
X_14115_ clknet_leaf_78_clk _01228_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08522__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ net2426 net177 net396 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
X_14046_ clknet_leaf_84_clk _01159_ net1270 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14009__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ net2571 net164 net402 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11656__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ cpu.IM0.address_IM\[31\] _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06916__A1 cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net2434 net171 net411 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13033__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ net972 cpu.RF0.registers\[1\]\[0\] net806 vssd1 vssd1 vccd1 vccd1 _02711_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14133__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__A2 _02160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07351_ net524 _02641_ _02607_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o21a_2
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire784_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07282_ cpu.RF0.registers\[17\]\[7\] net605 _02555_ _02560_ _02561_ vssd1 vssd1 vccd1
+ vccd1 _02573_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07644__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09021_ cpu.RF0.registers\[13\]\[31\] net659 _04303_ _04304_ _04306_ vssd1 vssd1
+ vccd1 vccd1 _04312_ sky130_fd_sc_hd__a2111o_1
XANTENNA_max_cap834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12516__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 cpu.FetchedInstr\[1\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 cpu.RF0.registers\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold223 cpu.DM0.readdata\[5\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 cpu.RF0.registers\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 a1.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 a1.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10036__A cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold267 cpu.RF0.registers\[17\]\[29\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 cpu.RF0.registers\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ cpu.IM0.address_IM\[7\] cpu.IM0.address_IM\[6\] _05189_ vssd1 vssd1 vccd1
+ vccd1 _05209_ sky130_fd_sc_hd__and3_1
XANTENNA__09825__A _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_6
Xhold289 cpu.RF0.registers\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout714 _02007_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08357__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_A _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_2
X_09854_ _04446_ _05142_ _05143_ cpu.CU0.funct3\[0\] cpu.CU0.funct3\[2\] vssd1 vssd1
+ vccd1 vccd1 _05145_ sky130_fd_sc_hd__a311o_1
Xfanout758 _02186_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1104_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_4
XANTENNA__12959__Q a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06887__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ net1083 cpu.RF0.registers\[22\]\[19\] net852 vssd1 vssd1 vccd1 vccd1 _04096_
+ sky130_fd_sc_hd__and3_1
X_09785_ _03634_ _04051_ _04053_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout564_A _05640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ net955 cpu.RF0.registers\[2\]\[23\] net769 vssd1 vssd1 vccd1 vccd1 _02288_
+ sky130_fd_sc_hd__and3_1
X_08736_ _03996_ _04026_ _03995_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_20_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_72_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S cpu.DM0.next_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ cpu.RF0.registers\[20\]\[2\] net709 net652 cpu.RF0.registers\[7\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ net1036 cpu.RF0.registers\[22\]\[13\] net800 vssd1 vssd1 vccd1 vccd1 _02909_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07883__A2 _02162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ cpu.RF0.registers\[23\]\[4\] _02045_ _03874_ _03875_ _03876_ vssd1 vssd1
+ vccd1 vccd1 _03889_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10219__A1 cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10219__B2 cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07511__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ net973 cpu.RF0.registers\[11\]\[8\] net777 vssd1 vssd1 vccd1 vccd1 _02840_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07096__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net1132 net1605 net912 _05667_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__a31o_1
XANTENNA__08832__B2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09219_ net453 _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__or2_1
X_10491_ net1483 net918 net750 a1.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 _00164_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12426__A cpu.DM0.data_i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ cpu.LCD0.row_1\[100\] _06024_ _06034_ cpu.LCD0.row_2\[28\] _06126_ vssd1
+ vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08596__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ cpu.LCD0.row_1\[121\] _06014_ _06051_ _06060_ _01961_ vssd1 vssd1 vccd1 vccd1
+ _06061_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_9_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ net2541 net219 net418 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
X_12092_ cpu.LCD0.nextState\[3\] cpu.LCD0.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _05993_
+ sky130_fd_sc_hd__and2_2
Xhold790 cpu.RF0.registers\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13056__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__B _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ net1924 net224 net429 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__mux2_1
XANTENNA__14301__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A0 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07255__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__A2 _04405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ clknet_leaf_22_clk net1528 net1172 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1490 cpu.RF0.registers\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net2896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__A2 _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__B2 a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14451__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ net2610 net173 net321 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14664_ cpu.LCD0.lcd_en vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08086__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net2451 net209 net326 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13615_ clknet_leaf_87_clk _00728_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08517__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net506 _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__and3_1
XANTENNA__07421__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14595_ clknet_leaf_61_clk _01697_ net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07087__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ clknet_leaf_102_clk _00659_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net990 _04774_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__nand2_1
XANTENNA__08373__X _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ clknet_leaf_95_clk _00590_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10689_ net2488 net2557 net902 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ cpu.DM0.data_i\[22\] net534 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08252__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12383__B2 cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ net1122 net1607 net531 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__a21o_1
XANTENNA__11386__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ clknet_leaf_104_clk _01142_ net1156 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_06920_ cpu.IG0.Instr\[27\] net634 net519 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a21o_1
XANTENNA__13549__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ net1038 cpu.RF0.registers\[24\]\[27\] net812 vssd1 vssd1 vccd1 vccd1 _02142_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _04807_ _04854_ _04860_ net278 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a22o_1
XANTENNA__09839__B1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06782_ cpu.RF0.registers\[9\]\[30\] net699 net651 cpu.RF0.registers\[7\]\[30\] _02018_
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08521_ net1106 cpu.RF0.registers\[25\]\[6\] net864 vssd1 vssd1 vccd1 vccd1 _03812_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10449__B2 a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13699__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12010__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ net1094 cpu.RF0.registers\[30\]\[8\] net839 vssd1 vssd1 vccd1 vccd1 _03743_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07865__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ cpu.RF0.registers\[13\]\[0\] net598 _02691_ _02692_ _02693_ vssd1 vssd1 vccd1
+ vccd1 _02694_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09067__A1 _04357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07331__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ net1093 cpu.RF0.registers\[27\]\[10\] net879 vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout145_A _05839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ net1063 cpu.RF0.registers\[30\]\[3\] net763 vssd1 vssd1 vccd1 vccd1 _02625_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ net980 cpu.RF0.registers\[10\]\[7\] net788 vssd1 vssd1 vccd1 vccd1 _02556_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08290__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_A _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ net934 cpu.RF0.registers\[5\]\[31\] net866 vssd1 vssd1 vccd1 vccd1 _04295_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07196_ net1051 cpu.RF0.registers\[27\]\[10\] net777 vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_83_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13079__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08162__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12374__B2 cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__Y _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12680__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07059__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14324__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1319_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout681_A _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
Xfanout511 net513 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11296__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__B net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ net625 _05073_ net1022 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__o21a_1
Xfanout522 net525 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_8
Xfanout533 _05848_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10053__X _05328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
Xfanout555 _01965_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07075__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _05126_ _05127_ _03079_ net443 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__o2bb2a_1
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14474__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout588 _02169_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_6
Xfanout599 _02154_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_8
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09768_ _05016_ _05030_ _05043_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09290__A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08719_ cpu.RF0.registers\[16\]\[0\] net635 _04007_ _04008_ _04009_ vssd1 vssd1 vccd1
+ vccd1 _04010_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07803__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ net438 _04358_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_1_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ cpu.RF0.registers\[21\]\[31\] net129 net346 vssd1 vssd1 vccd1 vccd1 _01143_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ net1956 net144 net357 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XANTENNA__07241__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__Q cpu.DM0.data_i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13400_ clknet_leaf_18_clk _00513_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net2477 net2263 net898 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
X_14380_ clknet_leaf_32_clk _01491_ net1245 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07608__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06706__X cpu.RU0.next_read_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ net2322 net161 net364 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_62_clk _00444_ net1309 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10543_ net47 net916 vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[1\] net1245 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10474_ net25 net755 _05640_ a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12365__B2 cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _06104_ _06110_ net556 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ clknet_leaf_35_clk _00373_ net1259 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08033__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ cpu.LCD0.row_2\[17\] _06003_ _06036_ cpu.LCD0.row_1\[17\] _06043_ vssd1 vssd1
+ vccd1 vccd1 _06044_ sky130_fd_sc_hd__a221o_1
XANTENNA__09781__A2 _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12075_ cpu.LCD0.cnt_500hz\[13\] cpu.LCD0.cnt_500hz\[12\] _05974_ vssd1 vssd1 vccd1
+ vccd1 _05978_ sky130_fd_sc_hd__and3_1
XANTENNA__10404__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__X _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net2002 net925 net273 _05903_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07416__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12977_ clknet_leaf_44_clk net1488 net1303 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09297__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ net2082 _05845_ net322 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07847__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13991__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14647_ clknet_leaf_22_clk _01748_ net1173 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07151__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ net2496 net145 net332 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ clknet_leaf_50_clk net2209 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_29 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13529_ clknet_leaf_92_clk _00642_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14347__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07050_ cpu.RF0.registers\[9\]\[19\] net573 _02319_ _02321_ _02324_ vssd1 vssd1 vccd1
+ vccd1 _02341_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_11_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XANTENNA__10367__B1 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13371__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14497__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12939__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ net1098 cpu.RF0.registers\[17\]\[29\] net884 vssd1 vssd1 vccd1 vccd1 _03243_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12005__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06511__B cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ net963 cpu.RF0.registers\[11\]\[27\] net776 vssd1 vssd1 vccd1 vccd1 _02194_
+ sky130_fd_sc_hd__and3_1
X_07883_ cpu.RF0.registers\[21\]\[29\] _02162_ net589 cpu.RF0.registers\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a22o_1
XANTENNA__07326__C net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ net495 _03233_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__nand2_1
X_06834_ _01848_ net633 _02123_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06846__D_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__X _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ net292 _04652_ _04657_ _04770_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__o211a_1
X_06765_ net938 net855 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08504_ _03783_ _03788_ _03792_ _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__nor4_1
XANTENNA__07299__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _03732_ _03769_ _04040_ _04045_ _03733_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a311o_2
XANTENNA__07838__A2 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ net36 net35 net38 net37 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__nor4_1
XFILLER_0_91_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ cpu.RF0.registers\[14\]\[9\] net650 _03724_ _03725_ net665 vssd1 vssd1 vccd1
+ vccd1 _03726_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07061__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ cpu.RF0.registers\[29\]\[11\] net672 _03638_ _03640_ _03647_ vssd1 vssd1
+ vccd1 vccd1 _03657_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07317_ net982 cpu.RF0.registers\[1\]\[3\] net807 vssd1 vssd1 vccd1 vccd1 _02608_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09269__B net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09460__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ cpu.RF0.registers\[8\]\[13\] net708 net646 cpu.RF0.registers\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07248_ _02535_ _02536_ _02537_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__or4_1
XANTENNA__13714__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout896_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _02465_ _02467_ _02469_ _02439_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__o31a_2
XFILLER_0_24_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10190_ _02004_ _05146_ _05449_ _05453_ _05451_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08620__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1306 net1313 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14236__RESET_B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1317 net1322 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__buf_2
XANTENNA__13864__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 _05938_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_8
Xfanout1328 net1331 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__buf_2
Xfanout341 _05936_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_4
Xfanout1339 net1342 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09572__X _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout363 _05930_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout374 _05927_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_8
XANTENNA__07236__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 _05925_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12900_ clknet_leaf_26_clk _00089_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11754__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _05922_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_6
X_13880_ clknet_leaf_18_clk _00993_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ clknet_leaf_41_clk _00050_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09279__A1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12283__B1 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12762_ net1477 net498 net279 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ clknet_leaf_47_clk _01603_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ net2300 net195 net347 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
XANTENNA__13043__Q cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ net2199 cpu.LCD0.row_2\[87\] net1001 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10894__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13244__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14432_ clknet_leaf_16_clk _01543_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_30_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11644_ net2086 net203 net355 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14363_ clknet_leaf_58_clk net1424 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10597__A0 cpu.LCD0.row_1\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08254__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11575_ net1987 net221 net364 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__mux2_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[21\] net1170 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ net1132 net1637 net912 _05650_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13394__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14294_ clknet_leaf_57_clk _01407_ net1367 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ clknet_leaf_21_clk _00425_ net1173 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10457_ net6 net753 net563 net2824 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__o22a_1
XANTENNA__10833__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08006__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10349__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09195__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ clknet_leaf_34_clk _00356_ net1250 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10388_ net1126 _01797_ net266 vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ net744 _05987_ _05993_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09923__A cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ cpu.LCD0.cnt_500hz\[7\] _05966_ net502 vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08714__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _02271_ _05847_ net283 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09642__B _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06550_ net308 net728 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06481_ cpu.f0.state\[8\] _01872_ cpu.f0.next_lcd_en vssd1 vssd1 vccd1 vccd1 _00024_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08493__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08220_ _03509_ _03510_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_60_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13737__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08151_ _03439_ _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06506__B cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ cpu.RF0.registers\[13\]\[14\] net598 net569 cpu.RF0.registers\[10\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
X_08082_ _02274_ _03147_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload47_A clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11839__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07033_ net964 cpu.RF0.registers\[4\]\[19\] net781 vssd1 vssd1 vccd1 vccd1 _02324_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_77_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12524__A cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13887__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08984_ cpu.IM0.address_IM\[26\] net551 _04273_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_
+ sky130_fd_sc_hd__a22o_4
XANTENNA__10044__A cpu.IM0.address_IM\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13117__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ _03222_ _03223_ _03224_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__or4_1
XANTENNA__11574__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07866_ cpu.RF0.registers\[22\]\[28\] net604 net587 cpu.RF0.registers\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a22o_1
X_09605_ net494 _04037_ _04882_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a31o_2
XFILLER_0_79_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06817_ cpu.CU0.opcode\[6\] _01850_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ net1031 cpu.RF0.registers\[31\]\[22\] net827 vssd1 vssd1 vccd1 vccd1 _03088_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_35_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13267__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net292 _04626_ _04632_ _04770_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__o211a_1
XANTENNA__14512__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__B1 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06748_ net940 net852 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10815__A1 cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ net471 _04650_ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10918__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06679_ a1.CPU_DAT_O\[15\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[15\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_47_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ net1079 cpu.RF0.registers\[30\]\[9\] net837 vssd1 vssd1 vccd1 vccd1 _03709_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08184__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _04687_ _04688_ net470 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__B2 _06332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08615__C _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__A0 cpu.f0.write_data\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08349_ net1088 cpu.RF0.registers\[26\]\[11\] net860 vssd1 vssd1 vccd1 vccd1 _03640_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09433__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1341_X net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11360_ net2400 net180 net391 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06798__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ net1020 net540 _05539_ cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__a31o_1
XANTENNA__11749__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ net1785 net169 net399 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__mux2_1
XANTENNA__12434__A cpu.DM0.data_i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13030_ clknet_leaf_61_clk _00002_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__09736__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ _05491_ _05492_ net309 vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_56_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12740__A1 cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_1
X_10173_ _05436_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_37_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1114 cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 net1127 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_2
Xfanout1136 net1143 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14042__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13038__Q cpu.LCD0.row_1\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _05832_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_1
Xfanout1158 net1167 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11484__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout171 _05817_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
XANTENNA__06970__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_2
Xfanout182 net184 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ clknet_leaf_88_clk _01045_ net1290 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout193 _05804_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XANTENNA__10503__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07263__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ clknet_leaf_82_clk _00976_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12814_ clknet_leaf_37_clk _00033_ net1258 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14192__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__A1 _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12256__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ clknet_leaf_94_clk _00907_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10806__B2 _05751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12745_ _01795_ _01871_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08094__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ net2605 net2220 net1005 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ clknet_leaf_39_clk _01526_ net1254 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11627_ net1715 net151 net359 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__mux2_1
XANTENNA__08227__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ clknet_leaf_27_clk _01459_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09918__A cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__A2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ net2788 net177 net368 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11659__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 cpu.RF0.registers\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ net1450 net916 net751 a1.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 _00182_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09637__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold619 cpu.RF0.registers\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ clknet_leaf_10_clk _01390_ net1166 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10990__A0 cpu.f0.write_data\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ net1814 net167 net375 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09188__B1 _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ clknet_leaf_45_clk _00408_ net1312 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07438__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ clknet_leaf_53_clk net1601 net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1308 cpu.RF0.registers\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1319 cpu.RF0.registers\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06961__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ cpu.RF0.registers\[20\]\[17\] net594 _02989_ _02998_ _03000_ vssd1 vssd1
+ vccd1 vccd1 _03011_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09360__B1 _04650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _02903_ _02940_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06602_ net1350 _01973_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__nand2_2
XANTENNA__12247__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07582_ net1046 cpu.RF0.registers\[18\]\[12\] net770 vssd1 vssd1 vccd1 vccd1 _02873_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09321_ _04608_ _04611_ _04477_ _04567_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_14_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06533_ cpu.f0.num\[15\] _01808_ cpu.f0.num\[20\] _01813_ _01902_ vssd1 vssd1 vccd1
+ vccd1 _01922_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08716__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09252_ net473 _04521_ _04485_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__o21ai_1
X_06464_ a1.curr_state\[0\] _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08203_ cpu.RF0.registers\[11\]\[21\] net690 net659 cpu.RF0.registers\[13\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a22o_1
X_09183_ _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06395_ cpu.f0.num\[20\] vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A _05786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07426__B1 _02682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ cpu.RF0.registers\[11\]\[23\] net690 _03411_ _03414_ _03419_ vssd1 vssd1
+ vccd1 vccd1 _03425_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09828__A _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11569__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__A1 cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ cpu.RF0.registers\[28\]\[25\] net705 net672 cpu.RF0.registers\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a22o_1
XANTENNA__09547__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1134_A _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10981__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ cpu.RF0.registers\[26\]\[23\] net599 _02279_ _02286_ _02292_ vssd1 vssd1
+ vccd1 vccd1 _02307_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14065__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout594_A _02160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1301_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ net1077 cpu.RF0.registers\[19\]\[26\] net835 vssd1 vssd1 vccd1 vccd1 _04258_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout859_A _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07354__Y _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ net957 cpu.RF0.registers\[12\]\[30\] net765 vssd1 vssd1 vccd1 vccd1 _03209_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08898_ cpu.RF0.registers\[9\]\[17\] net699 net670 cpu.RF0.registers\[22\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ cpu.RF0.registers\[15\]\[24\] _02167_ net568 cpu.RF0.registers\[25\]\[24\]
+ _03124_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a221o_1
XANTENNA__13902__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_X net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07514__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__B1 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10860_ net1620 net216 net430 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09519_ _02758_ _04698_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_45_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ net989 cpu.f0.data_adr\[22\] vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12530_ _06301_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08345__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12461_ cpu.f0.i\[3\] _06256_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_95_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ clknet_leaf_7_clk _01313_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ net1656 net212 net383 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
X_12392_ net2752 cpu.DM0.data_i\[2\] net733 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14408__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11479__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ clknet_leaf_69_clk _01244_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11343_ net2753 net224 net391 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ clknet_leaf_1_clk _01175_ net1142 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ net2401 net242 net400 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__mux2_1
X_13013_ clknet_leaf_36_clk _00202_ net1264 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10225_ cpu.f0.i\[6\] _05477_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a21o_1
XANTENNA__10724__A0 cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14558__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ cpu.IM0.address_IM\[26\] _05411_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 cpu.DM0.state\[1\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10412__A cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ cpu.IM0.address_IM\[20\] net931 _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _00043_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08089__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__X _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__B2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13582__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ clknet_leaf_13_clk _01028_ net1241 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09893__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08696__A2 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12229__B1 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13846_ clknet_leaf_58_clk _00959_ net1368 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13777_ clknet_leaf_76_clk _00890_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08448__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _02347_ net533 net283 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07656__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12728_ _01776_ cpu.DM0.dhit cpu.f0.state\[7\] net986 _01759_ vssd1 vssd1 vccd1 vccd1
+ _01720_ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07120__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12659_ cpu.LCD0.row_2\[61\] cpu.LCD0.row_2\[53\] net997 vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09948__A2 _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14088__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11389__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 cpu.RF0.registers\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ clknet_leaf_56_clk _01442_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold416 cpu.RF0.registers\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 a1.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 cpu.RF0.registers\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold449 cpu.RF0.registers\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout907 net911 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _02101_ _05043_ _05159_ _05160_ cpu.IM0.pc_enable vssd1 vssd1 vccd1 vccd1
+ _05161_ sky130_fd_sc_hd__o221a_1
Xfanout918 net924 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_2
Xfanout929 _00017_ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12180__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ cpu.RF0.registers\[31\]\[19\] net687 net651 cpu.RF0.registers\[7\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13925__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 cpu.RF0.registers\[12\]\[7\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 cpu.RF0.registers\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _03732_ _03769_ _03733_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1127 cpu.RF0.registers\[20\]\[29\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 cpu.LCD0.row_2\[81\] vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10322__A cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1149 cpu.LCD0.row_1\[48\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07703_ net959 cpu.RF0.registers\[1\]\[17\] net805 vssd1 vssd1 vccd1 vccd1 _02994_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08683_ cpu.RF0.registers\[1\]\[1\] net713 net669 cpu.RF0.registers\[22\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a22o_1
XANTENNA__07334__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08687__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07634_ net1045 cpu.RF0.registers\[18\]\[13\] net770 vssd1 vssd1 vccd1 vccd1 _02925_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10494__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__B _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07895__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07631__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ cpu.RF0.registers\[16\]\[8\] net581 _02835_ _02839_ _02842_ vssd1 vssd1 vccd1
+ vccd1 _02856_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout342_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ net484 net470 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__nand2_1
X_06516_ cpu.f0.num\[9\] _01799_ cpu.f0.num\[30\] _01821_ vssd1 vssd1 vccd1 vccd1
+ _01905_ sky130_fd_sc_hd__a2bb2o_1
X_07496_ cpu.RF0.registers\[10\]\[5\] net570 _02773_ _02775_ _02779_ vssd1 vssd1 vccd1
+ vccd1 _02787_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13305__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ _04524_ _04525_ net475 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06447_ net1411 _01780_ _01854_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10992__A _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__A _02865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09939__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ net464 _03766_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06378_ cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__inv_2
XANTENNA__08462__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11299__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08117_ net935 cpu.RF0.registers\[4\]\[23\] net874 vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ net465 _04276_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08048_ _03337_ _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
Xhold950 cpu.RF0.registers\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07509__C net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 cpu.RF0.registers\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 cpu.RF0.registers\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 cpu.LCD0.row_1\[43\] vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10931__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold994 cpu.RF0.registers\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12171__A2 _06019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ cpu.IM0.address_IM\[14\] net931 _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _00037_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09293__A _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09999_ _05276_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__B1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ cpu.RF0.registers\[28\]\[31\] net128 net318 vssd1 vssd1 vccd1 vccd1 _01367_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13316__Q cpu.DM0.data_i\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13700_ clknet_leaf_95_clk _00813_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10912_ cpu.DM0.readdata\[24\] _05107_ net739 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__mux2_1
X_14680_ net1402 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__10485__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net1718 net146 net329 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07350__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ clknet_leaf_0_clk _00744_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10843_ net2686 net243 net431 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13562_ clknet_leaf_93_clk _00675_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10774_ cpu.IM0.address_IM\[17\] net1013 net284 _05728_ vssd1 vssd1 vccd1 vccd1 _05729_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07102__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ cpu.f0.i\[21\] net1019 _06289_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and3_1
XANTENNA__14230__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ clknet_leaf_73_clk _00606_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ cpu.DM0.data_i\[30\] net535 vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08803__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ net1120 net1455 net529 cpu.IG0.Instr\[17\] vssd1 vssd1 vccd1 vccd1 _01501_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__B1 _05683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14380__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06604__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14114_ clknet_leaf_94_clk _01227_ net1227 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11326_ net2791 net152 net394 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11937__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ clknet_leaf_89_clk _01158_ net1280 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10841__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ net2279 net168 net403 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__mux2_1
XANTENNA__07169__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10208_ _02102_ net521 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__o21a_1
XANTENNA__07716__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ net2252 net187 net412 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__mux2_1
XANTENNA__06916__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12972__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ cpu.IM0.address_IM\[24\] _03143_ _05398_ vssd1 vssd1 vccd1 vccd1 _05407_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07154__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08669__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11672__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13328__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ clknet_leaf_8_clk _00942_ net1164 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10228__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11425__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07350_ cpu.RF0.registers\[0\]\[3\] net618 _02637_ _02640_ vssd1 vssd1 vccd1 vccd1
+ _02641_ sky130_fd_sc_hd__o22a_2
XFILLER_0_85_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07281_ cpu.RF0.registers\[8\]\[7\] net612 _02550_ _02551_ _02562_ vssd1 vssd1 vccd1
+ vccd1 _02572_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08841__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ cpu.RF0.registers\[14\]\[31\] net650 _04295_ _04300_ _04302_ vssd1 vssd1
+ vccd1 vccd1 _04311_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14102__RESET_B net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08282__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 cpu.RF0.registers\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12008__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold213 cpu.RF0.registers\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _01521_ vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 cpu.SR1.char_in\[0\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 cpu.RF0.registers\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold257 cpu.RF0.registers\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11847__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold268 cpu.RF0.registers\[25\]\[7\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net717 net135 _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold279 cpu.RF0.registers\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12532__A cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 _02020_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_2
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_2
XANTENNA__12153__A2 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07014__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout737 _01853_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_2
X_09853_ _04446_ _05142_ _05143_ _04449_ cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1
+ _05144_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_42_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07626__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__A1 cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06907__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 _02186_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08804_ cpu.RF0.registers\[6\]\[19\] net676 _04092_ _04093_ _04094_ vssd1 vssd1 vccd1
+ vccd1 _04095_ sky130_fd_sc_hd__a2111o_1
XANTENNA__14103__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _04863_ _04881_ _05074_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__or3_1
X_06996_ net955 cpu.RF0.registers\[11\]\[23\] net775 vssd1 vssd1 vccd1 vccd1 _02287_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08735_ net467 _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__or2_2
XANTENNA__07064__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1299_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08666_ cpu.RF0.registers\[11\]\[2\] net689 net655 cpu.RF0.registers\[2\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a22o_1
XANTENNA__10467__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08457__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14253__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07617_ net964 cpu.RF0.registers\[15\]\[13\] net827 vssd1 vssd1 vccd1 vccd1 _02908_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09609__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ cpu.RF0.registers\[3\]\[4\] net643 net635 cpu.RF0.registers\[16\]\[4\] _03887_
+ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout724_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ net973 cpu.RF0.registers\[9\]\[8\] net759 vssd1 vssd1 vccd1 vccd1 _02839_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07479_ net1060 cpu.RF0.registers\[18\]\[5\] net772 vssd1 vssd1 vccd1 vccd1 _02770_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10926__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1254_X net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09218_ net465 net445 _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__o21ai_1
X_10490_ net1541 net918 net750 a1.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 _00163_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08192__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12845__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ net456 _04439_ _04436_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07399__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ _06053_ _06055_ _06057_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07239__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11757__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ net1778 net221 net420 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XANTENNA__12995__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ cpu.LCD0.row_2\[88\] _05983_ _05986_ cpu.LCD0.row_1\[80\] _05991_ vssd1 vssd1
+ vccd1 vccd1 _05992_ sky130_fd_sc_hd__a221o_1
Xhold780 cpu.LCD0.row_2\[56\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06711__Y _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 cpu.RF0.registers\[26\]\[30\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12144__A2 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ net2632 net230 net429 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__mux2_1
XANTENNA__08899__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07571__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12993_ clknet_leaf_22_clk net1451 net1171 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11492__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1480 a1.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 net2886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1491 cpu.f0.data_adr\[23\] vssd1 vssd1 vccd1 vccd1 net2897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09312__A3 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ net2098 net195 net320 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14663_ net1387 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__07702__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ net1560 net204 net327 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__mux2_1
XANTENNA__12604__A0 cpu.LCD0.row_2\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13614_ clknet_leaf_2_clk _00727_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13620__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ cpu.IG0.Instr\[10\] cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__and2_2
X_14594_ clknet_leaf_52_clk _01696_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10757_ net2872 net561 net536 _05716_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__a22o_1
XANTENNA__10836__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13545_ clknet_leaf_106_clk _00658_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08823__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ clknet_leaf_98_clk _00589_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ cpu.LCD0.row_1\[94\] net2684 net908 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_91_clk_X clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13770__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ net1826 net731 net501 _06237_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ net1122 net1966 net531 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07149__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11667__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ net2725 net230 net396 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
XANTENNA__14126__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ cpu.LCD0.row_2\[15\] _05998_ _06025_ cpu.LCD0.row_1\[63\] _06182_ vssd1 vssd1
+ vccd1 vccd1 _06183_ sky130_fd_sc_hd__a221o_1
X_14028_ clknet_leaf_87_clk _01141_ net1287 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07446__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ net1053 net813 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13150__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14276__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ cpu.RF0.registers\[17\]\[30\] net694 _02032_ _02034_ _02043_ vssd1 vssd1
+ vccd1 vccd1 _02072_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09839__A1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ net949 cpu.RF0.registers\[12\]\[6\] net869 vssd1 vssd1 vccd1 vccd1 _03811_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08277__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07314__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ net945 cpu.RF0.registers\[7\]\[8\] net845 vssd1 vssd1 vccd1 vccd1 _03742_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_44_clk_X clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06509__B cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07402_ net1048 cpu.RF0.registers\[27\]\[0\] net777 vssd1 vssd1 vccd1 vccd1 _02693_
+ sky130_fd_sc_hd__and3_1
X_08382_ net1093 cpu.RF0.registers\[25\]\[10\] net863 vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12868__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ net1061 cpu.RF0.registers\[29\]\[3\] net793 vssd1 vssd1 vccd1 vccd1 _02624_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08724__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06825__A1 cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ net980 cpu.RF0.registers\[13\]\[7\] net794 vssd1 vssd1 vccd1 vccd1 _02555_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09003_ _03302_ _04289_ _04290_ _03271_ _03237_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__o311a_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_102_clk_X clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07195_ net1051 cpu.RF0.registers\[21\]\[10\] net797 vssd1 vssd1 vccd1 vccd1 _02486_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A cpu.IG0.Instr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _06230_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_2
XANTENNA__09527__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ net127 _05188_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__o21ai_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07356__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout523 net525 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_6
XANTENNA__14619__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout674_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_4
Xfanout556 _01961_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_4
X_09836_ _03080_ net434 _04923_ net293 net288 vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__o221a_1
XANTENNA__11885__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 _02193_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_8
Xfanout578 _02182_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_6
Xfanout589 _02169_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09767_ _05050_ _05051_ _05057_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__o21ai_4
X_06979_ _02259_ _02262_ _02264_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout841_A _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08718_ cpu.RF0.registers\[23\]\[0\] net1096 net845 vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13643__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09698_ _02213_ _04243_ _04915_ _04987_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o221a_1
XANTENNA__08187__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07305__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07091__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08618__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ net1104 cpu.RF0.registers\[25\]\[2\] net863 vssd1 vssd1 vccd1 vccd1 _03940_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14095__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07856__A3 _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ net1808 net149 net355 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XANTENNA__14024__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09058__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ net2288 cpu.LCD0.row_1\[25\] net908 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13793__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ net2105 net177 net364 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ clknet_leaf_61_clk _00443_ net1346 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ net1132 a1.ADR_I\[15\] net912 _05658_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08353__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14425__Q cpu.DM0.readdata\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13261_ clknet_leaf_33_clk cpu.RU0.next_FetchedInstr\[0\] net1246 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[0\] sky130_fd_sc_hd__dfrtp_1
X_10473_ net23 net753 net563 net2875 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__o22a_1
XANTENNA__14149__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ _05986_ _06106_ _06109_ _06075_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__or4b_1
XFILLER_0_32_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13192_ clknet_leaf_36_clk _00372_ net1264 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08650__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ cpu.LCD0.row_2\[105\] _06012_ _06031_ cpu.LCD0.row_1\[25\] vssd1 vssd1 vccd1
+ vccd1 _06043_ sky130_fd_sc_hd__a22o_1
XANTENNA__13173__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ cpu.LCD0.cnt_500hz\[12\] _05974_ cpu.LCD0.cnt_500hz\[13\] vssd1 vssd1 vccd1
+ vccd1 _05977_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11025_ cpu.f0.write_data\[30\] _05902_ net985 vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10420__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12976_ clknet_leaf_28_clk net1503 net1184 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
X_11927_ net2668 net136 net322 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
XANTENNA__07432__C net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14646_ clknet_leaf_21_clk _01747_ net1173 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11858_ net1525 net150 net331 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XANTENNA__08825__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ net287 _05752_ _05753_ net1016 cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1
+ vccd1 _05754_ sky130_fd_sc_hd__a32o_1
XANTENNA__08257__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_19 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ clknet_leaf_50_clk net2360 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ net2318 net177 net340 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13528_ clknet_leaf_7_clk _00641_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08009__B1 cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13459_ clknet_leaf_68_clk _00572_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__X _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__10367__A1 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13516__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07951_ net1099 cpu.RF0.registers\[27\]\[29\] net879 vssd1 vssd1 vccd1 vccd1 _03242_
+ sky130_fd_sc_hd__and3_1
X_06902_ net963 net776 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__inv_2
XANTENNA__07463__X _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ _01849_ _02085_ _02092_ net626 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__and4_1
X_09621_ net495 _03233_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__or2_1
X_09552_ net277 _04836_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a211o_1
XANTENNA__11619__A1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06764_ net936 cpu.RF0.registers\[13\]\[30\] net848 vssd1 vssd1 vccd1 vccd1 _02055_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12021__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08503_ cpu.RF0.registers\[17\]\[7\] net694 net673 cpu.RF0.registers\[29\]\[7\] _03793_
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ _04756_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08496__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06695_ a1.CPU_DAT_O\[31\] net889 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[31\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11860__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08434_ cpu.RF0.registers\[15\]\[9\] net682 _03704_ _03707_ _03709_ vssd1 vssd1 vccd1
+ vccd1 _03725_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ cpu.RF0.registers\[2\]\[11\] net656 _03637_ _03644_ _03646_ vssd1 vssd1 vccd1
+ vccd1 _03656_ sky130_fd_sc_hd__a2111o_1
XANTENNA__13046__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout422_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ net544 _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__or2_1
X_08296_ cpu.RF0.registers\[15\]\[13\] net682 net674 cpu.RF0.registers\[6\]\[13\]
+ _03578_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08173__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ cpu.RF0.registers\[8\]\[9\] net611 _02510_ _02527_ _02529_ vssd1 vssd1 vccd1
+ vccd1 _02538_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1331_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ _02458_ _02459_ _02460_ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout791_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08470__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14441__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A _01951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11100__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1307 net1309 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07517__C net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_8
Xfanout1318 net1322 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 _05938_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
Xfanout1329 net1331 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__clkbuf_4
Xfanout342 net345 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout353 _05933_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout364 _05930_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_8
Xfanout375 _05927_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09920__B1 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net389 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
X_09819_ net479 _04631_ _05040_ _04496_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__o211a_1
Xfanout397 _05922_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14205__RESET_B net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ clknet_leaf_14_clk _00049_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08348__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ cpu.f0.write_data\[19\] net497 net279 net1020 vssd1 vssd1 vccd1 vccd1 _01740_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11770__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ clknet_leaf_47_clk _01602_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11712_ net2653 net200 net346 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
X_12692_ net2452 cpu.LCD0.row_2\[86\] net1006 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XANTENNA__08645__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06717__X _02008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__B _04683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ net1997 net212 net355 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
X_14431_ clknet_leaf_17_clk _01542_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09436__C1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11574_ cpu.RF0.registers\[17\]\[7\] net226 net365 vssd1 vssd1 vccd1 vccd1 _00991_
+ sky130_fd_sc_hd__mux2_1
X_14362_ clknet_leaf_58_clk _01475_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13539__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13840__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
X_10525_ net69 net921 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13313_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[20\] net1169 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14293_ clknet_leaf_73_clk _01406_ net1341 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09476__A _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ clknet_leaf_22_clk _00424_ net1172 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ net5 net753 net563 net2886 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08380__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ clknet_leaf_37_clk _00355_ net1303 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10387_ net1127 _05611_ net266 net2799 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13689__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12126_ _05982_ _05989_ _05995_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__and3_4
XANTENNA__06973__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _05966_ net502 _05965_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__and3b_1
XANTENNA__09923__B cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ net1481 net926 net274 _05891_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a22o_1
XANTENNA__09415__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12959_ clknet_leaf_28_clk _00148_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13069__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11680__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__X _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14314__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06480_ cpu.K0.keyvalid _01870_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_83_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07686__D1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14629_ clknet_leaf_26_clk _01730_ net1182 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08150_ net445 _03437_ _03438_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__and3b_1
XANTENNA__14464__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07101_ _02386_ _02387_ _02391_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12906__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09386__A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ net1040 cpu.RF0.registers\[19\]\[19\] net821 vssd1 vssd1 vccd1 vccd1 _02323_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_77_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06803__A cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08721__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12016__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10325__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06522__B cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ cpu.RF0.registers\[0\]\[26\] net661 net547 vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10760__A1 _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__B2 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__Y _04683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ cpu.RF0.registers\[4\]\[30\] net586 _03201_ _03210_ _03217_ vssd1 vssd1 vccd1
+ vccd1 _03225_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07634__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07865_ cpu.RF0.registers\[17\]\[28\] net606 net595 cpu.RF0.registers\[7\]\[28\]
+ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__a221o_1
XANTENNA__10512__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _04477_ net272 _04884_ _04890_ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06816_ _02095_ _02090_ _02083_ cpu.CU0.opcode\[3\] vssd1 vssd1 vccd1 vccd1 _02107_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07796_ net1032 cpu.RF0.registers\[26\]\[22\] net786 vssd1 vssd1 vccd1 vccd1 _03087_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _04821_ _04825_ net479 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__mux2_1
X_06747_ net1117 net1110 net1112 net1115 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__and4bb_4
XANTENNA__12265__B2 cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07072__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11590__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ net472 _04721_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nand2_1
X_06678_ a1.CPU_DAT_O\[14\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10815__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12017__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08417_ cpu.RF0.registers\[10\]\[9\] net691 net638 cpu.RF0.registers\[26\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__a22o_1
XANTENNA__07800__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _04499_ _04501_ net453 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1167_X net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ net944 cpu.RF0.registers\[12\]\[11\] net868 vssd1 vssd1 vccd1 vccd1 _03639_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10579__A1 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10934__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ net1082 cpu.RF0.registers\[22\]\[13\] net851 vssd1 vssd1 vccd1 vccd1 _03570_
+ sky130_fd_sc_hd__and3_1
X_10310_ net540 _05549_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__nand2_1
XANTENNA__13831__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07995__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09296__A _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net2156 net181 net400 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _01801_ _05485_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07747__A2 _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10172_ cpu.IM0.address_IM\[28\] _03170_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10751__A1 _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1108 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11765__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12450__A cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1137 net1139 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout1148 net1211 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout161 _05832_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout1159 net1162 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_4
Xfanout172 _05817_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
XANTENNA__07544__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
X_13931_ clknet_leaf_90_clk _01044_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout194 _05804_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08172__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14337__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13862_ clknet_leaf_7_clk _00975_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12813_ clknet_leaf_37_clk _00032_ net1262 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ clknet_leaf_66_clk _00906_ net1293 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10806__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12744_ cpu.f0.write_data\[4\] net497 _01769_ _01770_ vssd1 vssd1 vccd1 vccd1 _01725_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07132__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13361__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__Q cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14487__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08806__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ cpu.LCD0.row_2\[77\] cpu.LCD0.row_2\[69\] net997 vssd1 vssd1 vccd1 vccd1
+ _01668_ sky130_fd_sc_hd__mux2_1
XANTENNA__07710__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ clknet_leaf_31_clk net1437 net1249 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ net2530 net157 net358 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14345_ clknet_leaf_27_clk _01458_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09918__B cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ net2482 net153 net366 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
XANTENNA__08632__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10508_ net94 net922 net747 net1412 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold609 cpu.RF0.registers\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
X_11488_ net2161 net183 net377 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
X_14276_ clknet_leaf_97_clk _01389_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10439_ net1125 _05637_ net264 net2120 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__a2bb2o_1
X_13227_ clknet_leaf_3_clk _00407_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12192__B1 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09493__X _04784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__A cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13158_ clknet_leaf_54_clk net1681 net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07157__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__A1 cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ _05981_ _05982_ net744 _06009_ cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1
+ _06010_ sky130_fd_sc_hd__a32o_1
X_13089_ clknet_leaf_48_clk _00269_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[53\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12360__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1309 cpu.LCD0.row_1\[16\] vssd1 vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06996__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__inv_2
XANTENNA__09360__B2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ cpu.LCD0.currentState\[1\] cpu.LCD0.nextState\[1\] net555 vssd1 vssd1 vccd1
+ vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07581_ net1046 cpu.RF0.registers\[31\]\[12\] _02129_ vssd1 vssd1 vccd1 vccd1 _02872_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09320_ _03118_ net434 net288 _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__o211a_1
X_06532_ _01809_ cpu.f0.i\[17\] _01815_ net1018 _01904_ vssd1 vssd1 vccd1 vccd1 _01921_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08285__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07123__B1 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ net296 _04541_ _04540_ _04539_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__o211a_1
X_06463_ a1.WRITE_I a1.READ_I vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14437__D net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ _03479_ _03490_ _03491_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09182_ _03964_ _03992_ net463 vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06394_ cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08133_ cpu.RF0.registers\[31\]\[23\] net687 _03409_ _03410_ _03416_ vssd1 vssd1
+ vccd1 vccd1 _03424_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07426__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__B _04813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ net943 cpu.RF0.registers\[2\]\[25\] net854 vssd1 vssd1 vccd1 vccd1 _03355_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07629__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10981__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07015_ cpu.RF0.registers\[4\]\[23\] net586 _02288_ _02290_ _02293_ vssd1 vssd1 vccd1
+ vccd1 _02306_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08451__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07067__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11585__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13234__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ net1080 cpu.RF0.registers\[23\]\[26\] net844 vssd1 vssd1 vccd1 vccd1 _04257_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12486__A1 cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ net1029 cpu.RF0.registers\[30\]\[30\] net762 vssd1 vssd1 vccd1 vccd1 _03208_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ _04184_ _04185_ _04186_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__or4_1
XANTENNA__08154__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10497__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ cpu.RF0.registers\[27\]\[24\] net592 net585 cpu.RF0.registers\[2\]\[24\]
+ _03125_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a221o_1
XANTENNA__07901__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10929__S net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ cpu.RF0.registers\[2\]\[21\] net584 _03052_ _03053_ _03059_ vssd1 vssd1 vccd1
+ vccd1 _03070_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_49_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09518_ _02758_ _04401_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10790_ net989 _04617_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__nand2_1
XANTENNA__08195__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09449_ _03335_ _03371_ _04275_ _04243_ net460 net452 vssd1 vssd1 vccd1 vccd1 _04740_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08862__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12460_ _06256_ _06257_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08923__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ net2773 net216 net382 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
X_12391_ cpu.DM0.readdata\[1\] cpu.DM0.data_i\[1\] net733 vssd1 vssd1 vccd1 vccd1
+ _01517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07968__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ net2887 net230 net391 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
X_14130_ clknet_leaf_60_clk _01243_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14433__Q cpu.DM0.readdata\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14061_ clknet_leaf_101_clk _01174_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11273_ net2075 net246 net400 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__mux2_1
XANTENNA__12174__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ clknet_leaf_28_clk _00201_ net1190 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
X_10224_ cpu.K0.keyvalid cpu.f0.state\[5\] _01870_ net728 vssd1 vssd1 vccd1 vccd1
+ _05479_ sky130_fd_sc_hd__a31o_2
XANTENNA__10724__A1 _05030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ cpu.IM0.address_IM\[26\] _05411_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__Q cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 a1.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13727__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ net626 _05096_ net1023 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__o21a_1
XANTENNA__07705__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10488__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ clknet_leaf_94_clk _01027_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09893__A2 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13845_ clknet_leaf_74_clk _00958_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10839__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13877__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13776_ clknet_leaf_75_clk _00889_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07105__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988_ net1425 net926 net274 _05877_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06459__A2 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ cpu.f0.state\[2\] cpu.f0.state\[7\] _06251_ vssd1 vssd1 vccd1 vccd1 _01759_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07440__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09929__A cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12658_ cpu.LCD0.row_2\[60\] cpu.LCD0.row_2\[52\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01651_ sky130_fd_sc_hd__mux2_1
XANTENNA__13107__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ net2422 net216 net358 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12589_ net721 net134 net932 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_74_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14328_ clknet_leaf_57_clk _01441_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold406 cpu.RF0.registers\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 a1.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 cpu.RF0.registers\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 cpu.RF0.registers\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ clknet_leaf_68_clk _01372_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12165__B1 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10715__A1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net911 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06919__B1 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout919 net924 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ cpu.RF0.registers\[28\]\[19\] net705 net666 vssd1 vssd1 vccd1 vccd1 _04111_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09383__B _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 cpu.LCD0.row_2\[43\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 cpu.RF0.registers\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__inv_2
XANTENNA__12468__A1 cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1128 cpu.RF0.registers\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07615__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10322__B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1139 cpu.RF0.registers\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14652__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10479__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07702_ net1028 cpu.RF0.registers\[30\]\[17\] net761 vssd1 vssd1 vccd1 vccd1 _02993_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ cpu.RF0.registers\[17\]\[1\] net695 net658 cpu.RF0.registers\[13\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07633_ net1037 cpu.RF0.registers\[26\]\[13\] net786 vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12089__X _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08727__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_A _05822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ cpu.RF0.registers\[22\]\[8\] net604 net595 cpu.RF0.registers\[7\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ net480 net474 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06515_ _01815_ net1018 cpu.f0.num\[24\] _01817_ vssd1 vssd1 vccd1 vccd1 _01904_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_17_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07495_ cpu.RF0.registers\[16\]\[5\] net582 _02764_ _02766_ _02772_ vssd1 vssd1 vccd1
+ vccd1 _02786_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12581__A1_N _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout335_A _05937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06446_ cpu.DM0.enable _01779_ _01851_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__or3b_1
XFILLER_0_5_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _04365_ _04418_ net451 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10992__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14032__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ _04454_ _04455_ net454 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
X_06377_ cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09558__B _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1244_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__inv_2
X_09096_ net465 _04243_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08047_ net446 _03336_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__X _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold940 cpu.RF0.registers\[31\]\[5\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12156__B1 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold951 cpu.RF0.registers\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 a1.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold973 cpu.RF0.registers\[19\]\[25\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 _00259_ vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 cpu.RF0.registers\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__A2 _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ cpu.IM0.address_IM\[14\] _02385_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12459__A1 cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ cpu.RF0.registers\[1\]\[27\] net714 _04237_ _04238_ _04239_ vssd1 vssd1 vccd1
+ vccd1 _04240_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__09324__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ net2224 net136 net318 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__mux2_1
X_10911_ net2115 net153 net430 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net2709 net150 net327 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13630_ clknet_leaf_86_clk _00743_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10842_ _05180_ _05777_ net721 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_15_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08356__C net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13561_ clknet_leaf_92_clk _00674_ net1239 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07260__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10773_ cpu.f0.data_adr\[17\] _04734_ net989 vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12512_ cpu.f0.i\[21\] _06289_ _06290_ net262 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__o211a_1
XANTENNA__09749__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08653__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ clknet_leaf_70_clk _00605_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06725__X _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12443_ cpu.DM0.readdata\[29\] net730 net500 _06245_ vssd1 vssd1 vccd1 vccd1 _01545_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14525__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ net1119 net2883 net530 cpu.IG0.Instr\[16\] vssd1 vssd1 vccd1 vccd1 _01500_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09260__B1 _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08091__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ clknet_leaf_64_clk _01226_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11325_ net2641 net165 net394 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12147__B1 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11256_ net2664 net184 net404 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__mux2_1
X_14044_ clknet_leaf_8_clk _01157_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10158__C1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08366__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ _05468_ _05469_ cpu.IM0.address_IM\[30\] net930 vssd1 vssd1 vccd1 vccd1 _00053_
+ sky130_fd_sc_hd__a2bb2o_1
X_11187_ cpu.RF0.registers\[5\]\[17\] net192 net410 vssd1 vssd1 vccd1 vccd1 _00617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ cpu.IM0.address_IM\[25\] _02272_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07435__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11953__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ _05341_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__nor2_1
X_13828_ clknet_leaf_96_clk _00941_ net1231 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14055__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13759_ clknet_leaf_0_clk _00872_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ cpu.RF0.registers\[23\]\[7\] net613 _02548_ _02549_ _02557_ vssd1 vssd1 vccd1
+ vccd1 _02571_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_73_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_X clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 cpu.RF0.registers\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 cpu.RF0.registers\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold225 cpu.RF0.registers\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 cpu.LCD0.row_1\[126\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold247 cpu.RF0.registers\[9\]\[8\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 cpu.RF0.registers\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _05205_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__xnor2_1
Xhold269 cpu.RF0.registers\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout705 _02017_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_6
XANTENNA__08357__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 net718 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_4
Xfanout727 _01938_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12024__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _04516_ _04684_ _04715_ _05141_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and4_1
Xfanout738 net740 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_2
X_08803_ net1083 cpu.RF0.registers\[25\]\[19\] net862 vssd1 vssd1 vccd1 vccd1 _04094_
+ sky130_fd_sc_hd__and3_1
X_09783_ _04896_ _05005_ _05059_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or4b_1
X_06995_ net955 cpu.RF0.registers\[13\]\[23\] net790 vssd1 vssd1 vccd1 vccd1 _02286_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout285_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08734_ cpu.IM0.address_IM\[0\] net553 _04023_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_59_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08665_ _03952_ _03953_ _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07616_ net1045 cpu.RF0.registers\[20\]\[13\] net781 vssd1 vssd1 vccd1 vccd1 _02907_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_49_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09609__A2 _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ cpu.RF0.registers\[10\]\[4\] net692 net681 cpu.RF0.registers\[18\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12613__A1 cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ net1052 cpu.RF0.registers\[19\]\[8\] net823 vssd1 vssd1 vccd1 vccd1 _02838_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout717_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14548__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07096__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ net981 cpu.RF0.registers\[8\]\[5\] net814 vssd1 vssd1 vccd1 vccd1 _02769_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09217_ net460 net446 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__or2_1
X_06429_ cpu.c0.count\[9\] cpu.c0.count\[10\] _01835_ vssd1 vssd1 vccd1 vccd1 _01840_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11103__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ _04437_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__nor2_1
XANTENNA__13572__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__B2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _04368_ _04369_ net455 vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11110_ net2847 net226 net421 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XANTENNA__09508__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12090_ cpu.LCD0.row_2\[64\] _05988_ _05990_ cpu.LCD0.row_2\[80\] vssd1 vssd1 vccd1
+ vccd1 _05991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 cpu.RF0.registers\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _01647_ vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 cpu.f0.num\[21\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net2435 net232 net429 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11352__A1 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07255__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13327__Q cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12992_ clknet_leaf_44_clk net1413 net1304 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A2 _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07552__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 cpu.LCD0.cnt_20ms\[1\] vssd1 vssd1 vccd1 vccd1 net2876 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1481 cpu.RF0.registers\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net2887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 cpu.RF0.registers\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net2898 sky130_fd_sc_hd__dlygate4sd3_1
X_11943_ net1689 net198 net318 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14662_ net72 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
X_11874_ net1571 net213 net329 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__mux2_1
XANTENNA__08086__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13613_ clknet_leaf_101_clk _00726_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ cpu.IG0.Instr\[7\] cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__and2_2
X_14593_ clknet_leaf_50_clk net2405 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_13544_ clknet_leaf_98_clk _00657_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07087__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ net284 _05714_ _05715_ net1017 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1
+ vccd1 _05716_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08383__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08814__C net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__A1 cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ clknet_leaf_79_clk _00588_ net1314 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10687_ cpu.LCD0.row_1\[93\] cpu.LCD0.row_1\[101\] net900 vssd1 vssd1 vccd1 vccd1
+ _00317_ sky130_fd_sc_hd__mux2_1
XANTENNA__10418__A cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11013__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ cpu.DM0.data_i\[21\] net535 vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11948__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ cpu.DM0.enable net1122 net736 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__nor3_1
X_11308_ net2756 net233 net397 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12288_ cpu.LCD0.row_2\[95\] _05983_ _06021_ cpu.LCD0.row_1\[95\] vssd1 vssd1 vccd1
+ vccd1 _06182_ sky130_fd_sc_hd__a22o_1
XANTENNA__14621__Q cpu.f0.write_data\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ clknet_leaf_91_clk _01140_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11239_ net2145 net247 net404 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__mux2_1
XANTENNA__07011__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11683__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06780_ cpu.RF0.registers\[11\]\[30\] net690 _02040_ net665 _02012_ vssd1 vssd1 vccd1
+ vccd1 _02071_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_26_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13445__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ net1094 cpu.RF0.registers\[28\]\[8\] net868 vssd1 vssd1 vccd1 vccd1 _03741_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07401_ net971 cpu.RF0.registers\[15\]\[0\] net830 vssd1 vssd1 vccd1 vccd1 _02692_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ net1093 cpu.RF0.registers\[21\]\[10\] net865 vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07332_ net1062 cpu.RF0.registers\[25\]\[3\] net759 vssd1 vssd1 vccd1 vccd1 _02623_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07078__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire887_A _02006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13595__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07263_ net1061 cpu.RF0.registers\[22\]\[7\] net802 vssd1 vssd1 vccd1 vccd1 _02554_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10328__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12019__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ _04287_ _04288_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07194_ net1051 cpu.RF0.registers\[20\]\[10\] net783 vssd1 vssd1 vccd1 vccd1 _02485_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10909__A1 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__S net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10762__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ _02004_ _05146_ _05191_ net625 vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__o31a_1
Xfanout502 _05958_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_2
Xfanout513 _02120_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_4
Xfanout524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_2
XANTENNA__07538__B1 _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 _05847_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_2
Xfanout546 _02124_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout557 _05997_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
X_09835_ net298 _04923_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__nand2_1
Xfanout568 _02191_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_8
XANTENNA__14220__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07075__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A _02050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _05052_ _05053_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ _02265_ _02266_ _02267_ _02268_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__or4_1
XANTENNA__08468__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08717_ cpu.RF0.registers\[29\]\[0\] net1096 net849 vssd1 vssd1 vccd1 vccd1 _04008_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07803__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ _02250_ _04275_ _04587_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__or3b_1
XANTENNA__08502__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14370__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07091__B _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ net949 cpu.RF0.registers\[15\]\[2\] net858 vssd1 vssd1 vccd1 vccd1 _03939_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12812__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _03866_ _03868_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10937__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_X net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12598__A0 cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ net2715 net2617 net909 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ net1664 net153 net362 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06716__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net46 net919 vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12962__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06856__B_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09215__A0 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ clknet_leaf_28_clk cpu.RU0.next_read_i net1190 vssd1 vssd1 vccd1 vccd1 a1.READ_I
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ net22 net752 net562 a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__o22a_1
XANTENNA__08931__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11022__A0 cpu.f0.write_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _06107_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__or2_1
XANTENNA__08569__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ clknet_leaf_34_clk _00371_ net1253 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ net1383 _06041_ _06042_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__and3_1
XANTENNA__07547__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13318__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14441__Q cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ cpu.LCD0.cnt_500hz\[12\] _05974_ _05976_ vssd1 vssd1 vccd1 vccd1 _01444_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ net509 net534 net282 vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12599__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__A _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__C net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ clknet_leaf_36_clk net1484 net1260 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07713__C net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11926_ net2101 net142 net323 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ clknet_leaf_16_clk _01746_ net1197 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_11857_ net1887 net155 net330 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XANTENNA__10847__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__A_N _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ net989 cpu.f0.data_adr\[27\] vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__or2_1
X_14576_ clknet_leaf_53_clk _01678_ net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_11788_ net2265 net154 net338 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13527_ clknet_leaf_64_clk _00640_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10739_ net286 _05702_ _05703_ net1014 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1
+ vccd1 _05704_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13458_ clknet_leaf_60_clk _00571_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08009__B2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11678__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ cpu.DM0.data_i\[13\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__12363__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13389_ clknet_leaf_103_clk _00502_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__06999__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14243__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07950_ net1098 cpu.RF0.registers\[30\]\[29\] net840 vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__and3_1
X_06901_ net1039 cpu.RF0.registers\[25\]\[27\] net757 vssd1 vssd1 vccd1 vccd1 _02192_
+ sky130_fd_sc_hd__and3_1
X_07881_ _03169_ _03171_ net522 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_4
X_09620_ _04907_ _04910_ net277 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__o21a_1
X_06832_ net741 _02091_ net629 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or3_2
XANTENNA__14393__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07940__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _04383_ _04655_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nor2_1
X_06763_ net940 net848 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__and2_4
XANTENNA__07623__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08502_ cpu.RF0.registers\[28\]\[7\] net706 net692 cpu.RF0.registers\[10\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a22o_1
X_09482_ net278 _04537_ _04764_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a211o_1
XANTENNA__07299__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06694_ a1.CPU_DAT_O\[30\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[30\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__08575__X _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07920__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08433_ cpu.RF0.registers\[8\]\[9\] net708 net651 cpu.RF0.registers\[7\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a22o_1
XANTENNA__12097__X _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__B _04025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12985__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A _05776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09445__A0 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08364_ cpu.RF0.registers\[1\]\[11\] net714 net701 cpu.RF0.registers\[9\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a22o_1
XANTENNA__09996__A1 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ cpu.IG0.Instr\[10\] net742 _02208_ net1066 vssd1 vssd1 vccd1 vccd1 _02606_
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ cpu.RF0.registers\[31\]\[13\] net687 _03583_ _03584_ _03585_ vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07246_ cpu.RF0.registers\[26\]\[9\] net599 _02515_ _02520_ _02531_ vssd1 vssd1 vccd1
+ vccd1 _02537_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11588__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ cpu.RF0.registers\[2\]\[11\] net584 net578 cpu.RF0.registers\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13610__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout310 _05943_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_6
Xfanout1308 net1309 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__clkbuf_4
Xfanout1319 net1322 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
Xfanout321 _05941_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_6
Xfanout332 _05938_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_8
Xfanout343 net345 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout354 _05932_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_6
Xfanout365 _05930_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_4
Xfanout376 _05927_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_6
X_09818_ net306 _05041_ _04480_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o21a_1
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09920__B2 cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _05921_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_90_clk_X clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ net484 _04821_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__or2_1
XANTENNA__13760__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10818__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12760_ cpu.f0.write_data\[18\] net498 net279 cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1
+ _01739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12283__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__A _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11711_ net2363 net208 net349 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ cpu.LCD0.row_2\[93\] cpu.LCD0.row_2\[85\] net997 vssd1 vssd1 vccd1 vccd1
+ _01684_ sky130_fd_sc_hd__mux2_1
XANTENNA__14245__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14116__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ clknet_leaf_17_clk _01541_ net1193 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11642_ net2486 net217 net354 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
XANTENNA__10046__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ clknet_leaf_72_clk _01474_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11573_ net2621 net230 net365 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07998__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_13312_ clknet_leaf_19_clk cpu.RU0.next_FetchedData\[19\] net1180 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[19\] sky130_fd_sc_hd__dfrtp_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ net1132 net1602 net912 _05649_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__a31o_1
XANTENNA__13140__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06733__X _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14292_ clknet_leaf_72_clk _01405_ net1340 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14266__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11498__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ clknet_leaf_34_clk _00423_ net1253 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10455_ net4 net753 net563 a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__o22a_1
XANTENNA__09476__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ clknet_leaf_35_clk _00354_ net1259 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10386_ cpu.f0.i\[5\] net270 vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__nand2_1
XANTENNA__07708__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ cpu.LCD0.row_1\[96\] _06024_ _06025_ cpu.LCD0.row_1\[56\] _06023_ vssd1 vssd1
+ vccd1 vccd1 _06026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13290__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ cpu.LCD0.cnt_500hz\[5\] cpu.LCD0.cnt_500hz\[4\] cpu.LCD0.cnt_500hz\[6\] _01955_
+ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ cpu.f0.write_data\[24\] _05890_ net995 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__mux2_1
XANTENNA__08714__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_X clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__C net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_X clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11961__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ clknet_leaf_28_clk _00147_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12274__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ net1727 net208 net325 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XANTENNA__10577__S net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12889_ clknet_leaf_30_clk _00020_ net1207 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ clknet_leaf_31_clk _01729_ net1202 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14609__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14559_ clknet_leaf_56_clk _01661_ net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13250__Q a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09089__D _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ cpu.RF0.registers\[18\]\[14\] net580 _02388_ _02389_ _02390_ vssd1 vssd1
+ vccd1 vccd1 _02391_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ cpu.IM0.address_IM\[25\] net552 _03369_ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07453__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ net1040 cpu.RF0.registers\[31\]\[19\] net827 vssd1 vssd1 vccd1 vccd1 _02322_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13633__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12734__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11201__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07187__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13550__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__C net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ _04262_ _04267_ _04271_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__or4_2
X_07933_ cpu.RF0.registers\[3\]\[30\] net609 _03204_ _03205_ _03208_ vssd1 vssd1 vccd1
+ vccd1 _03224_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07915__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13783__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__B cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10341__A cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07864_ cpu.RF0.registers\[2\]\[28\] net585 net577 cpu.RF0.registers\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09603_ _02830_ _03833_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06815_ _02102_ _02105_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_30_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ net959 cpu.RF0.registers\[15\]\[22\] net826 vssd1 vssd1 vccd1 vccd1 _03086_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout365_A _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14139__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _04823_ _04824_ net476 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__mux2_1
X_06746_ net944 net875 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__and2_2
XANTENNA__12265__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07650__A _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _03599_ _03600_ _04754_ _04755_ net493 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__o311a_1
X_06677_ a1.CPU_DAT_O\[13\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[13\]
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1274_A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08416_ net935 cpu.RF0.registers\[1\]\[9\] net882 vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13163__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09396_ _04455_ _04498_ net454 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08347_ net1088 cpu.RF0.registers\[20\]\[11\] net874 vssd1 vssd1 vccd1 vccd1 _03638_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08278_ cpu.RF0.registers\[5\]\[13\] net702 net671 cpu.RF0.registers\[23\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07229_ net1035 cpu.RF0.registers\[27\]\[9\] net775 vssd1 vssd1 vccd1 vccd1 _02520_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11111__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07097__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10240_ _01801_ _05485_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08944__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ cpu.IM0.address_IM\[28\] _03170_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_2
Xfanout1116 cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 cpu.f0.state\[6\] vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
Xfanout140 _05841_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__B cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout151 _05837_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08157__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_4
Xfanout162 _05832_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dlymetal6s2s_1
X_13930_ clknet_leaf_101_clk _01043_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10251__A cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout173 net176 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
Xfanout184 _05819_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10503__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 _05804_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ clknet_leaf_10_clk _00974_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07263__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11781__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ clknet_leaf_37_clk _00031_ net1262 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_100_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12256__A2 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13792_ clknet_leaf_9_clk _00905_ net1160 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06728__X _02019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08656__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _06342_ _01763_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12674_ cpu.LCD0.row_2\[76\] cpu.LCD0.row_2\[68\] net1002 vssd1 vssd1 vccd1 vccd1
+ _01667_ sky130_fd_sc_hd__mux2_1
XANTENNA__07683__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14413_ clknet_leaf_32_clk _01524_ net1254 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08094__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ net2667 net159 net358 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13656__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ clknet_leaf_27_clk _01457_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09487__A _04399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ net1784 net166 net366 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10975__C1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ net1479 net920 net749 a1.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 _00180_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ clknet_leaf_77_clk _01388_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10426__A cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ net2326 net172 net375 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XANTENNA__09188__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_104_clk _00406_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10438_ cpu.f0.i\[31\] net268 vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__nand2_1
XANTENNA__07438__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11956__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ clknet_leaf_51_clk _00337_ net1379 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10860__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10369_ net1127 cpu.f0.state\[5\] vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10742__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net744 _05993_ _05996_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__and3_4
X_13088_ clknet_leaf_48_clk _00268_ net1361 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[52\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ cpu.LCD0.cnt_20ms\[15\] cpu.LCD0.cnt_20ms\[14\] _05953_ _05954_ vssd1 vssd1
+ vccd1 vccd1 _05955_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10161__A cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09950__A cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13245__Q a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14167__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ cpu.LCD0.nextState\[0\] cpu.LCD0.currentState\[0\] net556 vssd1 vssd1 vccd1
+ vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XANTENNA__12247__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07580_ net1045 cpu.RF0.registers\[22\]\[12\] net801 vssd1 vssd1 vccd1 vccd1 _02871_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13186__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06531_ cpu.f0.num\[4\] _01794_ _01820_ cpu.f0.i\[30\] _01905_ vssd1 vssd1 vccd1
+ vccd1 _01920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _03195_ net448 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__xor2_1
X_06462_ net1 net915 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08201_ cpu.RF0.registers\[12\]\[21\] net696 net674 cpu.RF0.registers\[6\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__a22o_1
X_09181_ net469 _03992_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nor2_1
X_06393_ cpu.f0.i\[17\] vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14581__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ cpu.RF0.registers\[19\]\[23\] net640 _03412_ _03413_ _03418_ vssd1 vssd1
+ vccd1 vccd1 _03423_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07426__A2 _02716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09820__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload52_A clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__C _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ net1092 cpu.RF0.registers\[30\]\[25\] net839 vssd1 vssd1 vccd1 vccd1 _03354_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12027__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07014_ cpu.RF0.registers\[6\]\[23\] net583 _02280_ _02298_ net621 vssd1 vssd1 vccd1
+ vccd1 _02305_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10055__B _05328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1022_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ net934 cpu.RF0.registers\[12\]\[26\] net867 vssd1 vssd1 vccd1 vccd1 _04256_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07916_ net1030 cpu.RF0.registers\[23\]\[30\] net816 vssd1 vssd1 vccd1 vccd1 _03207_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08896_ cpu.RF0.registers\[13\]\[17\] net659 net651 cpu.RF0.registers\[7\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__a22o_1
XANTENNA__07347__D1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__A cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__CLK clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ cpu.RF0.registers\[21\]\[24\] net593 net577 cpu.RF0.registers\[28\]\[24\]
+ _03126_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12238__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08476__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ cpu.RF0.registers\[10\]\[21\] net569 _03051_ _03062_ _03065_ vssd1 vssd1
+ vccd1 vccd1 _03069_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_49_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06729_ net943 net865 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07811__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_A _01860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11106__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ _04737_ _04738_ net476 vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09379_ _04668_ _04669_ net455 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11749__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11410_ net2273 net220 net385 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12390_ net1536 cpu.DM0.data_i\[0\] net733 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__mux2_1
XANTENNA__12410__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11341_ net2231 net234 net391 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13401__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14060_ clknet_leaf_87_clk _01173_ net1287 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ net2172 net251 net401 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ clknet_leaf_28_clk _00200_ net1190 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13059__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ net1442 net728 _05478_ cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__a22o_1
XANTENNA__12461__A cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09246__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ net717 net134 _05419_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__a211oi_1
XANTENNA__14607__RESET_B net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 _00181_ vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net126 _05357_ _05354_ net628 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a211o_1
XANTENNA__09878__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14454__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13913_ clknet_leaf_42_clk _01026_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14260__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07353__A1 cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__B2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13844_ clknet_leaf_71_clk _00957_ net1340 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12229__A2 _05988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13775_ clknet_leaf_80_clk _00888_ net1285 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ cpu.f0.write_data\[18\] _05876_ net995 vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__mux2_1
XANTENNA__08302__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ net1561 net726 _00020_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06803__D_N cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12657_ net2338 cpu.LCD0.row_2\[51\] net998 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__mux2_1
XANTENNA__10855__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ net2023 net220 net361 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06634__A a1.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ cpu.IM0.address_IM\[0\] _02682_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09010__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__C net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14327_ clknet_leaf_57_clk _01440_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11539_ cpu.RF0.registers\[16\]\[5\] net233 net369 vssd1 vssd1 vccd1 vccd1 _00957_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10156__A cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 cpu.RF0.registers\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 cpu.RF0.registers\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09945__A cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold429 cpu.f0.num\[22\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ clknet_leaf_59_clk _01371_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11686__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ clknet_leaf_12_clk _00389_ net1223 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09664__B _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14189_ clknet_leaf_103_clk _01302_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 net911 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 cpu.LCD0.row_2\[96\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ _03699_ _03700_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__or2_1
XANTENNA__07184__B net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1118 cpu.LCD0.row_2\[65\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 cpu.RF0.registers\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ net954 cpu.RF0.registers\[13\]\[17\] net790 vssd1 vssd1 vccd1 vccd1 _02992_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08681_ cpu.RF0.registers\[9\]\[1\] net701 net698 cpu.RF0.registers\[12\]\[1\] _03969_
+ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08541__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ net960 cpu.RF0.registers\[8\]\[13\] net811 vssd1 vssd1 vccd1 vccd1 _02923_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13821__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07895__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08727__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ cpu.RF0.registers\[17\]\[8\] net605 _02834_ _02836_ _02838_ vssd1 vssd1 vccd1
+ vccd1 _02854_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07631__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ _04426_ _04434_ net475 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_1
X_06514_ cpu.f0.num\[31\] cpu.f0.i\[31\] vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07494_ cpu.RF0.registers\[17\]\[5\] net606 _02769_ _02770_ _02771_ vssd1 vssd1 vccd1
+ vccd1 _02785_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07647__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _04366_ _04368_ net455 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__mux2_1
X_06445_ net1118 cpu.CU0.opcode\[4\] cpu.CU0.opcode\[6\] _01847_ vssd1 vssd1 vccd1
+ vccd1 _01853_ sky130_fd_sc_hd__or4_1
XANTENNA__13971__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ _03534_ net442 net461 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__mux2_1
X_06376_ cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08462__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08072__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13201__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ net446 _03371_ net466 vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
XANTENNA__14327__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1237_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ net446 _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06831__X _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 cpu.LCD0.row_1\[14\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11596__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 cpu.RF0.registers\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 cpu.LCD0.row_1\[34\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 cpu.RF0.registers\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 cpu.RF0.registers\[30\]\[7\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 cpu.RF0.registers\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold996 cpu.LCD0.row_1\[111\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14477__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ cpu.IM0.address_IM\[14\] _02385_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__nand2_1
XANTENNA__07806__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ cpu.RF0.registers\[30\]\[27\] net660 net636 cpu.RF0.registers\[16\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ net1077 cpu.RF0.registers\[24\]\[17\] net870 vssd1 vssd1 vccd1 vccd1 _04170_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_99_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08532__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _05389_ _05826_ net719 vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__mux2_2
X_11890_ net2332 net155 net326 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__mux2_1
XANTENNA__07886__A2 _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ cpu.DM0.readdata\[4\] _05016_ net739 vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13560_ clknet_leaf_7_clk _00673_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10772_ a1.ADR_I\[16\] net558 net536 _05727_ vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07638__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08934__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ _05556_ _06267_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13491_ clknet_leaf_68_clk _00604_ net1323 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09101__Y _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12442_ cpu.DM0.data_i\[29\] net535 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14444__Q cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ net1123 net2044 net531 cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1 _01499_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09260__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10945__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ clknet_leaf_4_clk _01225_ net1159 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11324_ net1693 net169 net395 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
X_14043_ clknet_leaf_94_clk _01156_ net1227 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11255_ net1856 net170 net403 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ net630 _04516_ net932 vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ net2915 net205 net410 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__mux2_1
XANTENNA__07574__A1 _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10137_ cpu.IM0.address_IM\[25\] _02272_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13844__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ cpu.IM0.address_IM\[18\] _05319_ cpu.IM0.address_IM\[19\] vssd1 vssd1 vccd1
+ vccd1 _05342_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07451__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ clknet_leaf_79_clk _00940_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13994__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ clknet_leaf_85_clk _00871_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06916__X _02207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ cpu.LCD0.row_2\[111\] net1897 net1001 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__mux2_1
X_13689_ clknet_leaf_65_clk _00802_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06364__A cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10157__Y _05424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08282__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12386__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12386__B2 cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold204 cpu.RF0.registers\[29\]\[27\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 cpu.RF0.registers\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
X_14679__1401 vssd1 vssd1 vccd1 vccd1 _14679__1401/HI net1401 sky130_fd_sc_hd__conb_1
XANTENNA__13374__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 cpu.RF0.registers\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _00342_ vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09920_ _05183_ _05195_ _05196_ _02797_ cpu.IM0.address_IM\[6\] vssd1 vssd1 vccd1
+ vccd1 _05206_ sky130_fd_sc_hd__a32o_1
XANTENNA__11269__X _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 cpu.FetchedInstr\[24\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 cpu.RF0.registers\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06370__Y _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout706 _02017_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XANTENNA__07195__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 net718 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_4
X_09851_ _04551_ _04577_ _04601_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nor3b_1
Xfanout728 _01937_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07626__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout739 net740 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload15_A clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ net1083 cpu.RF0.registers\[17\]\[19\] net883 vssd1 vssd1 vccd1 vccd1 _04093_
+ sky130_fd_sc_hd__and3_1
X_09782_ net513 _05061_ _05066_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__o211a_2
XANTENNA__14111__RESET_B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ net1028 cpu.RF0.registers\[17\]\[23\] net804 vssd1 vssd1 vccd1 vccd1 _02285_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07923__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ cpu.RF0.registers\[0\]\[0\] net664 net549 vssd1 vssd1 vccd1 vccd1 _04024_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout180_A _05829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ cpu.RF0.registers\[30\]\[2\] _02053_ net644 cpu.RF0.registers\[3\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a22o_1
XANTENNA__10321__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07615_ net1036 cpu.RF0.registers\[17\]\[13\] net804 vssd1 vssd1 vccd1 vccd1 _02906_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08457__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07361__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ _03873_ _03884_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout445_A _03436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1187_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ net970 cpu.RF0.registers\[3\]\[8\] net823 vssd1 vssd1 vccd1 vccd1 _02837_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08754__A _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout612_A _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ net1061 cpu.RF0.registers\[20\]\[5\] net782 vssd1 vssd1 vccd1 vccd1 _02768_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08293__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09216_ net449 _04506_ _04505_ net301 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a211o_1
X_06428_ cpu.c0.count\[10\] _01837_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08192__C net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13717__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__B2 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ net463 _03931_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nor2_1
XANTENNA__12563__X _06329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06359_ net1453 vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_32_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09585__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ _03402_ net445 net466 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08029_ cpu.RF0.registers\[12\]\[24\] net698 net669 cpu.RF0.registers\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a22o_1
Xhold760 cpu.RF0.registers\[11\]\[17\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 cpu.RF0.registers\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 cpu.RF0.registers\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net2688 net243 net428 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
Xhold793 cpu.LCD0.row_2\[95\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ clknet_leaf_36_clk net1480 net1264 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
Xhold1460 cpu.K0.code\[6\] vssd1 vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08505__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1471 cpu.RF0.registers\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net2877 sky130_fd_sc_hd__dlygate4sd3_1
X_11942_ net1904 net210 net318 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
Xhold1482 cpu.RF0.registers\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net2888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07859__A2 _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1493 a1.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net2899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14661_ net72 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14439__Q cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ cpu.RF0.registers\[26\]\[9\] net216 net326 vssd1 vssd1 vccd1 vccd1 _01281_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07271__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13343__Q cpu.RF0.registers\[0\]\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13247__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06531__A2 _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ clknet_leaf_79_clk _00725_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10824_ cpu.IG0.Instr\[11\] _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__and2_1
X_14592_ clknet_leaf_53_clk _01694_ net1363 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ clknet_leaf_81_clk _00656_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ net990 cpu.f0.data_adr\[12\] vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09481__A1 _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__A2 _03042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13474_ clknet_leaf_10_clk _00587_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10686_ cpu.LCD0.row_1\[92\] cpu.LCD0.row_1\[100\] net903 vssd1 vssd1 vccd1 vccd1
+ _00316_ sky130_fd_sc_hd__mux2_1
XANTENNA__13397__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12368__B2 cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14642__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12425_ cpu.DM0.readdata\[20\] net730 net501 _06236_ vssd1 vssd1 vccd1 vccd1 _01536_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08036__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10715__B1_N net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09495__A _02473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ net2593 _06219_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__xor2_1
X_11307_ net2745 net243 net396 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
X_12287_ cpu.LCD0.row_2\[87\] _05990_ _06007_ cpu.LCD0.row_2\[119\] _06180_ vssd1
+ vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a221o_1
XANTENNA__09782__X _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ clknet_leaf_101_clk _01139_ net1213 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11238_ net2891 net251 net405 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__mux2_1
XANTENNA__07446__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ net503 _05910_ _05915_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and3_4
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07400_ net971 cpu.RF0.registers\[12\]\[0\] net767 vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14172__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08380_ net945 cpu.RF0.registers\[15\]\[10\] net857 vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_58_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07331_ net1061 cpu.RF0.registers\[22\]\[3\] net802 vssd1 vssd1 vccd1 vccd1 _02622_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07262_ net982 cpu.RF0.registers\[11\]\[7\] net777 vssd1 vssd1 vccd1 vccd1 _02553_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12359__A1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09001_ _03270_ _04290_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07193_ net1046 cpu.RF0.registers\[24\]\[10\] net812 vssd1 vssd1 vccd1 vccd1 _02484_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07918__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08983__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _05189_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nor2_1
XANTENNA__09527__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout503 _05909_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07356__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout525 _02125_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_4
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout536 net539 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
XANTENNA__12531__A1 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
XFILLER_0_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09834_ _04526_ net272 _04566_ _04532_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a22o_1
Xfanout558 net561 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1102_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _02190_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_6
X_09765_ _04535_ _04903_ _04998_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06977_ cpu.RF0.registers\[20\]\[25\] net594 net580 cpu.RF0.registers\[18\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
X_08716_ cpu.RF0.registers\[24\]\[0\] net1096 net871 vssd1 vssd1 vccd1 vccd1 _04007_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09696_ _03145_ net446 _04647_ _03371_ _02274_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o32a_1
XFILLER_0_83_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08187__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ cpu.RF0.registers\[8\]\[2\] net707 _03935_ _03936_ _03937_ vssd1 vssd1 vccd1
+ vccd1 _03938_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_1_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ _03866_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08484__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10058__C1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07529_ cpu.RF0.registers\[16\]\[6\] net582 _02801_ _02813_ _02817_ vssd1 vssd1 vccd1
+ vccd1 _02820_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08266__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11114__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ net1134 net2755 net914 _05657_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09215__A1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ net21 net752 net562 net1594 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ _06003_ _06027_ _06028_ _06034_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__or4_1
XANTENNA__07387__X _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13190_ clknet_leaf_34_clk _00370_ net1246 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06732__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12770__A1 cpu.f0.write_data\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net119 _01965_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__or2_1
XANTENNA__08974__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__B2 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10254__A cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10781__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ cpu.LCD0.cnt_500hz\[12\] _05974_ net502 vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a21boi_1
Xhold590 cpu.RF0.registers\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07266__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net1412 net926 net274 _05901_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14195__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ clknet_leaf_35_clk net1542 net1260 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12286__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1290 cpu.LCD0.row_1\[86\] vssd1 vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_2_clk_X clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ net2550 net144 net324 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XANTENNA__06504__A2 cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14678__1400 vssd1 vssd1 vccd1 vccd1 _14678__1400/HI net1400 sky130_fd_sc_hd__conb_1
X_14644_ clknet_leaf_24_clk _01745_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_11856_ net2674 net161 net331 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__mux2_1
XANTENNA__12589__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ net991 _04601_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nand2_1
XANTENNA__08825__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14575_ clknet_leaf_56_clk _01677_ net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08257__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11787_ net1863 net164 net338 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10738_ net987 cpu.f0.data_adr\[7\] vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__or2_2
XANTENNA__07465__B1 _02755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13526_ clknet_leaf_57_clk _00639_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11959__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_77_clk _00570_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10716__X _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ net2549 net1819 net898 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12408_ net1472 net732 _06227_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_11_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11013__A1 _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06642__A a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13388_ clknet_leaf_88_clk _00501_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14632__Q cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12761__A1 cpu.f0.write_data\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_12339_ net1423 _06208_ _06210_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11694__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ net1049 net759 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__and2_2
X_14009_ clknet_leaf_91_clk _01122_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09672__B _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13412__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _03170_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__inv_2
XANTENNA__14538__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__B1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ net514 net512 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__or2_4
XFILLER_0_78_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07940__A1 cpu.CU0.bit30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ net291 _04837_ _04840_ net298 _04839_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06762_ net1092 net839 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__and2_4
XFILLER_0_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08501_ _03775_ _03789_ _03790_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13562__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _02940_ _04766_ _04771_ net302 _04769_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o221ai_1
XANTENNA__08496__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06693_ a1.CPU_DAT_O\[29\] net889 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08432_ _03708_ _03720_ _03721_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__or4_1
XANTENNA_clkload82_A clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ cpu.RF0.registers\[15\]\[11\] net682 net674 cpu.RF0.registers\[6\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09445__A1 _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout143_A _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07314_ net524 _02602_ _02603_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__o21a_1
XANTENNA__11252__A1 _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ cpu.RF0.registers\[30\]\[13\] net660 _03574_ _03576_ _03577_ vssd1 vssd1
+ vccd1 vccd1 _03585_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11869__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ cpu.RF0.registers\[6\]\[9\] net583 _02512_ _02523_ _02525_ vssd1 vssd1 vccd1
+ vccd1 _02536_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_27_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout310_A _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12201__B1 _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ cpu.RF0.registers\[15\]\[11\] net590 _02466_ net621 vssd1 vssd1 vccd1 vccd1
+ _02467_ sky130_fd_sc_hd__a211o_1
XANTENNA__14068__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06552__A cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08470__C net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10763__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1317_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 _03564_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_4
XFILLER_0_26_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout311 _05943_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13092__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08708__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1309 net1313 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_2
Xfanout322 net325 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_6
Xfanout333 _05938_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_4
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_4
XANTENNA__08479__A _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 _05932_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout366 _05929_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09817_ _04198_ _04664_ _04200_ _04091_ _04208_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__o2111a_1
Xfanout377 _05927_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13905__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_6
XANTENNA__10521__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _05921_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10530__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12268__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ net483 _04825_ _05038_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10818__A1 cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09679_ _02604_ _03899_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ net1861 net202 net348 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10294__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ cpu.LCD0.row_2\[92\] cpu.LCD0.row_2\[84\] net1004 vssd1 vssd1 vccd1 vccd1
+ _01683_ sky130_fd_sc_hd__mux2_1
XANTENNA__12448__B cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09103__A _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ net1746 net221 net357 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__mux2_1
XANTENNA__09436__A1 _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__B2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ clknet_leaf_71_clk net1447 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11572_ net2898 net233 net365 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ clknet_leaf_20_clk cpu.RU0.next_FetchedData\[18\] net1176 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[18\] sky130_fd_sc_hd__dfrtp_1
X_10523_ net68 net918 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__and2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_14291_ clknet_leaf_68_clk _01404_ net1324 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12464__A cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ clknet_leaf_37_clk _00422_ net1306 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ net3 net755 _05640_ a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__a22o_1
XANTENNA__08947__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08380__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14452__Q cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ clknet_leaf_35_clk _00353_ net1261 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10385_ net1124 _05610_ net267 net2920 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13435__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12124_ _05984_ net743 _05987_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06973__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ cpu.LCD0.cnt_500hz\[5\] cpu.LCD0.cnt_500hz\[4\] _01955_ cpu.LCD0.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a31o_1
XANTENNA__08389__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _03142_ net533 net283 vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_70_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13585__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11019__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10809__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__B2 cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07135__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ clknet_leaf_21_clk _00146_ net1171 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11908_ net1564 net203 net324 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06637__A a1.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12888_ clknet_leaf_30_clk _00019_ net1202 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_83_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08555__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ clknet_leaf_31_clk _01728_ net1206 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ net2024 net222 net332 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__mux2_1
XANTENNA__11830__X _05938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14558_ clknet_leaf_47_clk _01660_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[69\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14210__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11689__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ clknet_leaf_3_clk _00622_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09667__B _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14489_ clknet_leaf_34_clk _01591_ net1253 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10993__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07030_ net964 cpu.RF0.registers\[13\]\[19\] net792 vssd1 vssd1 vccd1 vccd1 _02321_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12734__A1 _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08938__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12734__B2 cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__B1 _05688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14360__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ cpu.RF0.registers\[24\]\[26\] net684 net677 cpu.RF0.registers\[4\]\[26\]
+ _04250_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a221o_1
XANTENNA__13928__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06964__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ cpu.RF0.registers\[2\]\[30\] net584 _03200_ _03206_ _03215_ vssd1 vssd1 vccd1
+ vccd1 _03223_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12540__C cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ cpu.RF0.registers\[18\]\[28\] net579 net575 cpu.RF0.registers\[14\]\[28\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07634__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09602_ _02830_ _04402_ net291 _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a211o_1
X_06814_ _01850_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ net1032 cpu.RF0.registers\[17\]\[22\] net804 vssd1 vssd1 vccd1 vccd1 _03085_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ _04736_ _04795_ net457 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06745_ net1090 net855 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout358_A _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _03633_ _04051_ _03601_ _03632_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a211o_1
X_06676_ a1.CPU_DAT_O\[12\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_94_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13308__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__C net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ net1079 cpu.RF0.registers\[23\]\[9\] net844 vssd1 vssd1 vccd1 vccd1 _03706_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09395_ net512 _04289_ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_47_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1267_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08346_ net941 cpu.RF0.registers\[11\]\[11\] net880 vssd1 vssd1 vccd1 vccd1 _03637_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ net300 _03566_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__xor2_2
XANTENNA__09577__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07649__Y _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__C_N net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07228_ net959 cpu.RF0.registers\[11\]\[9\] net775 vssd1 vssd1 vccd1 vccd1 _02519_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07809__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07159_ net966 cpu.RF0.registers\[3\]\[11\] net821 vssd1 vssd1 vccd1 vccd1 _02450_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_56_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10170_ cpu.IM0.address_IM\[27\] net932 _05434_ _05435_ vssd1 vssd1 vccd1 vccd1 _00050_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_2
Xfanout1117 cpu.IG0.Instr\[15\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_1
XANTENNA__12489__B1 cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 _05845_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1139 net1143 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_2
Xfanout141 _05841_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_1
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout163 net166 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout174 net176 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07544__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _05804_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlymetal6s2s_1
X_13860_ clknet_leaf_99_clk _00973_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07380__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ clknet_leaf_37_clk _00030_ net1264 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10678__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ clknet_leaf_106_clk _00904_ net1136 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09104__Y _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12742_ _01794_ _01871_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07132__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14233__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12673_ net1755 net2399 net998 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XANTENNA__09409__A1 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__Q cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09409__B2 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14412_ clknet_leaf_37_clk _01523_ net1260 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10019__A2 _05140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ net2164 net178 net360 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XANTENNA__09768__A _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14343_ clknet_leaf_27_clk _01456_ net1184 vssd1 vssd1 vccd1 vccd1 cpu.K0.code\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ net2775 net169 net367 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__mux2_1
XANTENNA__08093__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire542 _03852_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08632__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14383__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ net1633 net916 net751 a1.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 _00179_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07840__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14274_ clknet_leaf_94_clk _01387_ net1222 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11486_ net1965 net185 net376 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__12825__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ clknet_leaf_74_clk _00405_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ _01820_ net268 _05636_ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10727__A0 cpu.f0.data_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ clknet_leaf_50_clk net1583 net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10368_ net526 _05594_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_72_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06946__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ cpu.LCD0.row_1\[32\] _06006_ _06007_ cpu.LCD0.row_2\[112\] _06005_ vssd1
+ vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__a221o_1
X_13087_ clknet_leaf_46_clk _00267_ net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ net541 _05539_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nand2_1
XANTENNA__09008__A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ cpu.LCD0.cnt_20ms\[17\] cpu.LCD0.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1 _05954_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11972__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06919__X _02210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13989_ clknet_leaf_103_clk _01102_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06530_ _01796_ cpu.f0.i\[6\] _01819_ cpu.f0.i\[29\] _01906_ vssd1 vssd1 vccd1 vccd1
+ _01919_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06367__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07123__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08285__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06461_ a1.curr_state\[2\] a1.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08200_ cpu.RF0.registers\[18\]\[21\] net680 net650 cpu.RF0.registers\[14\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13600__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11207__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ net469 _04025_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06392_ cpu.f0.num\[17\] vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__X _04321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ cpu.RF0.registers\[23\]\[23\] net671 _03408_ _03415_ _03417_ vssd1 vssd1
+ vccd1 vccd1 _03422_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06373__Y _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09820__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11212__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07198__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ net943 cpu.RF0.registers\[15\]\[25\] net857 vssd1 vssd1 vccd1 vccd1 _03353_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07831__B1 _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload45_A clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07013_ _02300_ _02301_ _02302_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__or4_1
XANTENNA__13750__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10194__A1 cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ net1077 cpu.RF0.registers\[28\]\[26\] net867 vssd1 vssd1 vccd1 vccd1 _04255_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1015_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ net1029 cpu.RF0.registers\[29\]\[30\] net791 vssd1 vssd1 vccd1 vccd1 _03206_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07364__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08895_ cpu.RF0.registers\[20\]\[17\] net710 net674 cpu.RF0.registers\[6\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12486__A3 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__B _02644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ cpu.RF0.registers\[20\]\[24\] _02160_ _03136_ net622 vssd1 vssd1 vccd1 vccd1
+ _03137_ sky130_fd_sc_hd__a211o_1
XANTENNA__07898__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07661__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14256__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ cpu.RF0.registers\[27\]\[21\] net591 _03048_ _03055_ _03056_ vssd1 vssd1
+ vccd1 vccd1 _03068_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout642_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1384_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08476__B _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09516_ net292 _04409_ net303 vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06728_ net1115 net1111 net1113 net1116 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08195__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09447_ _03402_ _03436_ _03471_ net443 net462 net455 vssd1 vssd1 vccd1 vccd1 _04738_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06659_ net1594 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[27\] sky130_fd_sc_hd__and2_1
XFILLER_0_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_clk_X clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13280__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09378_ _03471_ net440 net466 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12848__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08923__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ cpu.RF0.registers\[20\]\[12\] net710 _03607_ _03608_ _03610_ vssd1 vssd1
+ vccd1 vccd1 _03620_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_95_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08075__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09811__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11122__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11340_ net2230 net242 net391 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09100__B _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_X clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11271_ net2154 net253 net401 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__mux2_1
XANTENNA__12742__A _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_X clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ clknet_leaf_36_clk _00199_ net1263 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
X_10222_ cpu.f0.data_adr\[6\] net729 _05478_ cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1
+ _00059_ sky130_fd_sc_hd__a22o_1
XANTENNA__12174__A2 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _05416_ _05418_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nor2_1
XANTENNA__10262__A cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__B1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A gpio_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _05355_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__nor2_1
XANTENNA__09878__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 cpu.RF0.registers\[0\]\[10\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
X_13912_ clknet_leaf_6_clk _01025_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10488__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__X _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13843_ clknet_leaf_67_clk _00956_ net1298 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13623__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10986_ _02381_ net533 net282 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__o21ba_1
X_13774_ clknet_leaf_1_clk _00887_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07105__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12725_ net1529 cpu.LCD0.row_2\[119\] net1006 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08853__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ net2585 net2502 net999 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__mux2_1
XANTENNA__13773__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07289__Y _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ net2384 net225 net360 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
X_12587_ _06347_ net1789 _06320_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08605__A2 _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06634__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14326_ clknet_leaf_57_clk _01439_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11538_ net2491 net242 net368 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
XANTENNA__07449__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold408 cpu.RF0.registers\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11967__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold419 a1.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14129__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14257_ clknet_leaf_76_clk _01370_ net1335 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11469_ net2704 net254 net377 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12165__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ clknet_leaf_13_clk _00388_ net1237 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_14188_ clknet_leaf_88_clk _01301_ net1296 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13139_ clknet_leaf_53_clk _00319_ net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10172__A cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 cpu.RF0.registers\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 _01656_ vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ net1031 cpu.RF0.registers\[19\]\[17\] net820 vssd1 vssd1 vccd1 vccd1 _02991_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10479__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ net1103 cpu.RF0.registers\[20\]\[1\] net875 vssd1 vssd1 vccd1 vccd1 _03971_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07344__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ net959 cpu.RF0.registers\[11\]\[13\] net775 vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07912__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11207__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07562_ net1052 cpu.RF0.registers\[31\]\[8\] net830 vssd1 vssd1 vccd1 vccd1 _02853_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ net480 _04590_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__o21ai_1
X_06513_ cpu.f0.num\[26\] cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_17_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07493_ cpu.RF0.registers\[12\]\[5\] net571 _02763_ _02768_ _02777_ vssd1 vssd1 vccd1
+ vccd1 _02784_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_17_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09232_ net301 _04409_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06444_ net1118 cpu.CU0.opcode\[4\] cpu.CU0.opcode\[6\] _01847_ vssd1 vssd1 vccd1
+ vccd1 _01852_ sky130_fd_sc_hd__nor4_2
XFILLER_0_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09201__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _03629_ _03664_ net461 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__mux2_1
X_06375_ cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10347__A cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08114_ _03402_ _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nand2_1
X_09094_ net480 net475 vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07359__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11877__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ _03123_ _03145_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__xnor2_1
Xhold920 cpu.RF0.registers\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 _00238_ vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12156__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold942 cpu.RF0.registers\[21\]\[20\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 cpu.LCD0.row_2\[88\] vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 cpu.LCD0.row_1\[56\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__A1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 cpu.RF0.registers\[26\]\[8\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 cpu.LCD0.row_2\[33\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold997 _00335_ vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ cpu.IM0.address_IM\[13\] net931 _05274_ _05275_ vssd1 vssd1 vccd1 vccd1 _00036_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ cpu.RF0.registers\[12\]\[27\] net696 net690 cpu.RF0.registers\[11\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13646__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08878_ net1077 cpu.RF0.registers\[17\]\[17\] net882 vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08487__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ _02946_ _03021_ _03081_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__nor4_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11419__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net2315 net247 net432 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08218__B1_N net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13796__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09589__Y _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ net284 _05725_ _05726_ net1013 cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1
+ vccd1 _05727_ sky130_fd_sc_hd__a32o_1
XANTENNA__08296__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12510_ _05550_ _06268_ _06288_ net262 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__o211a_1
X_13490_ clknet_leaf_60_clk _00603_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09111__A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08653__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ cpu.DM0.readdata\[28\] net730 net500 _06244_ vssd1 vssd1 vccd1 vccd1 _01544_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13026__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12372_ net1122 net1457 net531 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 _01498_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07269__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14111_ clknet_leaf_106_clk _01224_ net1141 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11323_ net2612 net182 net397 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
XANTENNA__11787__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12147__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13176__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14042_ clknet_leaf_90_clk _01155_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11254_ net2013 net185 net404 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__mux2_1
XANTENNA__10158__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ net125 _05463_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a21oi_1
X_11185_ net2854 net173 net413 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10136_ _05403_ _05404_ cpu.IM0.address_IM\[24\] net932 vssd1 vssd1 vccd1 vccd1 _00047_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06782__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ cpu.IM0.address_IM\[19\] cpu.IM0.address_IM\[18\] _05319_ vssd1 vssd1 vccd1
+ vccd1 _05341_ sky130_fd_sc_hd__and3_1
XANTENNA__14571__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload1_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13826_ clknet_leaf_94_clk _00939_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13757_ clknet_leaf_66_clk _00870_ net1282 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10969_ net985 cpu.f0.write_data\[13\] vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10094__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ net2266 cpu.LCD0.row_2\[102\] net1006 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06645__A a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13688_ clknet_leaf_7_clk _00801_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14635__Q cpu.f0.write_data\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ net2499 net2392 net1009 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09787__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13519__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14309_ clknet_leaf_11_clk _01422_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold205 cpu.RF0.registers\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__B _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold216 a1.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold227 net92 vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 cpu.RF0.registers\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 cpu.RF0.registers\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06380__A cpu.f0.i\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14370__Q cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09850_ _05118_ _05121_ _05131_ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and4bb_1
XANTENNA__08211__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13669__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 _02014_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_8
Xfanout718 _02005_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_2
Xfanout729 _01937_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_0_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07565__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ net942 cpu.RF0.registers\[4\]\[19\] net875 vssd1 vssd1 vccd1 vccd1 _04092_
+ sky130_fd_sc_hd__and3_1
X_09781_ _04536_ _04564_ _04695_ _05071_ _05069_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a221oi_1
XPHY_EDGE_ROW_37_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06993_ net1027 cpu.RF0.registers\[28\]\[23\] net765 vssd1 vssd1 vccd1 vccd1 _02284_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10901__Y _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08732_ _04001_ _04006_ _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08663_ cpu.RF0.registers\[14\]\[2\] net649 net668 vssd1 vssd1 vccd1 vccd1 _03954_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10321__A1 cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14151__RESET_B net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07614_ net1045 cpu.RF0.registers\[23\]\[13\] net817 vssd1 vssd1 vccd1 vccd1 _02905_
+ sky130_fd_sc_hd__and3_1
X_08594_ cpu.RF0.registers\[14\]\[4\] net649 _03871_ _03877_ _03882_ vssd1 vssd1 vccd1
+ vccd1 _03885_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07545_ net973 cpu.RF0.registers\[14\]\[8\] net763 vssd1 vssd1 vccd1 vccd1 _02836_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10776__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout340_A _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ net1057 cpu.RF0.registers\[24\]\[5\] net813 vssd1 vssd1 vccd1 vccd1 _02767_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_46_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12276__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06427_ _01834_ _01836_ _01838_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[9\] sky130_fd_sc_hd__and3_1
X_09215_ net447 _04243_ net460 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_A _02144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ net467 _03964_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__nor2_1
X_06358_ cpu.f0.state\[2\] vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__inv_2
XANTENNA__13199__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14444__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07253__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ net444 net443 net466 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11400__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08028_ net1097 cpu.RF0.registers\[25\]\[24\] net863 vssd1 vssd1 vccd1 vccd1 _03319_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 cpu.RF0.registers\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 cpu.RF0.registers\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 cpu.LCD0.row_1\[15\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06721__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold783 cpu.RF0.registers\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _01686_ vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1302_X net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14594__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ cpu.IM0.address_IM\[10\] _02474_ _05247_ _05248_ vssd1 vssd1 vccd1 vccd1
+ _05260_ sky130_fd_sc_hd__a31oi_2
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ clknet_leaf_21_clk net1634 net1171 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1450 cpu.RF0.registers\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09106__A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1461 cpu.RF0.registers\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net2867 sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ cpu.RF0.registers\[28\]\[11\] net201 net319 vssd1 vssd1 vccd1 vccd1 _01347_
+ sky130_fd_sc_hd__mux2_1
Xhold1472 cpu.RF0.registers\[0\]\[1\] vssd1 vssd1 vccd1 vccd1 net2878 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__A1 cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1483 cpu.RF0.registers\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net2889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1494 cpu.LCD0.row_1\[105\] vssd1 vssd1 vccd1 vccd1 net2900 sky130_fd_sc_hd__dlygate4sd3_1
X_14660_ net72 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
X_11872_ net2381 net222 net329 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__mux2_1
X_13611_ clknet_leaf_90_clk _00724_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10686__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _02103_ _02123_ _02314_ net737 cpu.DM0.enable vssd1 vssd1 vccd1 vccd1 _05763_
+ sky130_fd_sc_hd__o32a_2
XANTENNA__08269__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14591_ clknet_leaf_55_clk net2447 net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08808__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12467__A cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13542_ clknet_leaf_7_clk _00655_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ net990 _04813_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nand2_1
XANTENNA__08009__X _03300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08383__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10685_ net2660 cpu.LCD0.row_1\[99\] net898 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
X_13473_ clknet_leaf_63_clk _00586_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12424_ cpu.DM0.data_i\[20\] net534 vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09495__B _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ _06219_ _06220_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11310__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13811__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11306_ net2738 net245 net397 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__mux2_1
X_12286_ cpu.LCD0.row_2\[127\] _06022_ _06030_ cpu.LCD0.row_1\[47\] vssd1 vssd1 vccd1
+ vccd1 _06180_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_73_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14025_ clknet_leaf_2_clk _01138_ net1154 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237_ net2628 net255 net405 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__mux2_1
X_11168_ net2586 net128 net414 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__mux2_1
XANTENNA__13961__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _05387_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__nor2_1
X_11099_ net2076 net142 net423 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__mux2_1
XANTENNA__08558__C net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11980__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14317__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07180__B1 _02004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12577__A2_N _06337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ clknet_leaf_77_clk _00922_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09457__C1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ net982 cpu.RF0.registers\[3\]\[3\] net823 vssd1 vssd1 vccd1 vccd1 _02621_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06375__A cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13341__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14467__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07261_ net1060 cpu.RF0.registers\[29\]\[7\] net793 vssd1 vssd1 vccd1 vccd1 _02552_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12909__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ _03271_ _03302_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07192_ net970 cpu.RF0.registers\[2\]\[10\] net771 vssd1 vssd1 vccd1 vccd1 _02483_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08590__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13491__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11220__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08983__A1 cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ cpu.IM0.address_IM\[5\] _05178_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout504 _05909_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_2
Xfanout526 _01893_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
X_09833_ net486 _04758_ _05062_ _04496_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__o211a_1
Xfanout548 _02087_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net458 net436 net290 _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__o211a_1
XANTENNA__10360__A cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06976_ cpu.RF0.registers\[19\]\[25\] net615 net572 cpu.RF0.registers\[12\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a22o_1
XANTENNA__08468__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08715_ _04002_ _04003_ _04004_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__or4_1
XANTENNA__07372__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09695_ _03172_ net447 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nor2_1
XANTENNA__11890__S net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_A _01965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ net1102 cpu.RF0.registers\[23\]\[2\] net846 vssd1 vssd1 vccd1 vccd1 _03937_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ _02795_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout722_A _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ cpu.RF0.registers\[19\]\[6\] net615 _02808_ _02811_ _02815_ vssd1 vssd1 vccd1
+ vccd1 _02819_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ cpu.RF0.registers\[29\]\[1\] net601 _02722_ _02726_ _02740_ vssd1 vssd1 vccd1
+ vccd1 _02750_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_92_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13834__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ net20 net754 net564 a1.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08931__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09129_ net467 _03766_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__nor2_1
XANTENNA__11130__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06732__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12140_ _05992_ _06002_ _06008_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or4_1
XANTENNA__10230__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07547__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10781__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13984__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ cpu.LCD0.cnt_500hz\[11\] _05973_ _05975_ net502 vssd1 vssd1 vccd1 vccd1 _01443_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 cpu.RF0.registers\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07529__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 cpu.RF0.registers\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ cpu.f0.write_data\[29\] _05900_ net995 vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13214__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10270__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ clknet_leaf_43_clk net1495 net1304 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13354__Q cpu.RF0.registers\[0\]\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1280 cpu.RF0.registers\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 cpu.RF0.registers\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
X_11924_ net1575 net150 net325 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06747__X _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13364__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14643_ clknet_leaf_23_clk _01744_ net1179 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11855_ net2169 net179 net332 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__mux2_1
XANTENNA__11305__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ a1.ADR_I\[26\] net558 net536 _05751_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__a22o_1
X_14574_ clknet_leaf_47_clk _01676_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[85\]
+ sky130_fd_sc_hd__dfstp_1
X_11786_ net1880 net167 net339 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__mux2_1
XANTENNA__07465__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13525_ clknet_leaf_68_clk _00638_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ net994 _04880_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__nand2_1
XANTENNA__08662__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ clknet_leaf_74_clk _00569_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10668_ net2316 cpu.LCD0.row_1\[82\] net902 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__mux2_1
XANTENNA__06923__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ cpu.DM0.data_i\[12\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10599_ cpu.LCD0.row_1\[5\] cpu.LCD0.row_1\[13\] net896 vssd1 vssd1 vccd1 vccd1 _00229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13387_ clknet_leaf_86_clk _00500_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06642__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12338_ cpu.LCD0.cnt_20ms\[12\] _06208_ net1369 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10772__A1 a1.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__B1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11975__S net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ cpu.LCD0.row_2\[86\] _05990_ _06019_ cpu.LCD0.row_1\[54\] vssd1 vssd1 vccd1
+ vccd1 _06164_ sky130_fd_sc_hd__a22o_1
X_14008_ clknet_leaf_6_clk _01121_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09390__A1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ net514 net512 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nor2_1
XANTENNA__10180__A _05443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07940__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13707__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ net1117 net1111 net1113 net1115 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__and4b_4
XANTENNA__07192__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10288__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ cpu.RF0.registers\[15\]\[7\] net683 net655 cpu.RF0.registers\[2\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09480_ net292 _04544_ _04770_ _04523_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__o211a_1
X_06692_ a1.CPU_DAT_O\[28\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08585__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ cpu.RF0.registers\[4\]\[9\] net677 _03705_ _03710_ _03714_ vssd1 vssd1 vccd1
+ vccd1 _03722_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07920__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08362_ cpu.RF0.registers\[18\]\[11\] net680 net636 cpu.RF0.registers\[16\]\[11\]
+ _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a221o_1
XANTENNA__13857__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07313_ net524 _02602_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_15_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload75_A clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ cpu.RF0.registers\[7\]\[13\] net651 _03572_ _03573_ net665 vssd1 vssd1 vccd1
+ vccd1 _03584_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07244_ cpu.RF0.registers\[25\]\[9\] net568 _02513_ _02519_ _02530_ vssd1 vssd1 vccd1
+ vccd1 _02535_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10460__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12881__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07175_ net1043 cpu.RF0.registers\[31\]\[11\] net830 net567 cpu.RF0.registers\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_41_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10355__A cpu.f0.i\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06552__B cpu.f0.state\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14584__RESET_B net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__A2 _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__C net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A1 cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11885__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13237__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _02759_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
Xfanout312 _05943_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_8
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout334 _05937_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A _02042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _05935_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout367 _05929_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_4
X_09816_ _04641_ _05097_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__o21bai_4
XANTENNA_hold1418_A a1.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 net381 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
Xfanout389 _05924_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_4
XANTENNA__07931__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__CLK clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _04384_ _04887_ _05037_ _04696_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14632__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ net543 _02248_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10818__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ net306 _03899_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08926__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ cpu.RF0.registers\[4\]\[3\] net678 net641 cpu.RF0.registers\[19\]\[3\] _03919_
+ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a221o_1
XANTENNA__08892__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11125__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11640_ net2244 net225 net356 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09436__A2 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ net2853 net241 net364 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07998__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13310_ clknet_leaf_19_clk cpu.RU0.next_FetchedData\[17\] net1176 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[17\] sky130_fd_sc_hd__dfrtp_1
X_10522_ net1132 net1622 net912 _05648_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__a31o_1
X_14290_ clknet_leaf_60_clk _01403_ net1344 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06743__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14012__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__B cpu.f0.i\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10453_ net33 net753 net563 net2930 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__o22a_1
X_13241_ clknet_leaf_26_clk _00421_ net1181 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10265__A cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06462__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13172_ clknet_leaf_36_clk _00352_ net1264 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10384_ cpu.f0.i\[4\] net271 vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07277__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11795__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ net743 _05989_ _05993_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12054_ _01961_ _05957_ _05964_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09372__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ net1977 net925 net273 _05889_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_70_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12956_ clknet_leaf_21_clk _00145_ net1171 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11907_ net1595 net213 net324 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12887_ clknet_leaf_28_clk _00018_ net1189 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06637__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14626_ clknet_leaf_30_clk _01727_ net1209 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11838_ net1674 net226 net333 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14557_ clknet_leaf_47_clk _01659_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08635__B1 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ net2734 net241 net340 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13508_ clknet_leaf_96_clk _00621_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_14488_ clknet_leaf_30_clk cpu.f0.next_write_i net1207 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_i
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10993__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ clknet_leaf_0_clk _00552_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14505__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12195__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07187__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__A1 cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__B _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ _04259_ _04268_ _04269_ _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07931_ cpu.RF0.registers\[27\]\[30\] net591 _03203_ _03209_ _03214_ vssd1 vssd1
+ vccd1 vccd1 _03222_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07915__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14655__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ cpu.RF0.registers\[19\]\[28\] net615 net601 cpu.RF0.registers\[29\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a22o_1
XANTENNA__08867__X _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09601_ net295 net299 _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06813_ _01778_ net1118 _01846_ _02083_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__o211a_1
X_07793_ net960 cpu.RF0.registers\[3\]\[22\] net820 vssd1 vssd1 vccd1 vccd1 _03084_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ _04796_ _04822_ net457 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06744_ net1116 net1110 net1112 net1114 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_17_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06828__A _02112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09463_ _03633_ _04051_ _03632_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a21oi_1
X_06675_ a1.CPU_DAT_O\[11\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[11\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ net1078 cpu.RF0.registers\[18\]\[9\] net855 vssd1 vssd1 vccd1 vccd1 _03705_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09394_ _03304_ _04287_ _04288_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and3_1
XANTENNA__14035__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07429__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ net1087 cpu.RF0.registers\[24\]\[11\] net870 vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08626__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout420_A _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1162_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08276_ net300 _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1270_A cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ net1036 cpu.RF0.registers\[19\]\[9\] net820 vssd1 vssd1 vccd1 vccd1 _02518_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14185__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07158_ net1043 cpu.RF0.registers\[29\]\[11\] net792 vssd1 vssd1 vccd1 vccd1 _02449_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07097__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_clk_X clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ _02369_ _02370_ _02371_ _02372_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__or4_1
XANTENNA__07394__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_2
Xfanout1129 cpu.f0.state\[4\] vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
Xfanout131 _05845_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
XANTENNA__08157__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 _05841_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_2
Xfanout186 _05814_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07904__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout197 net200 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
X_12810_ clknet_leaf_37_clk _00029_ net1266 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_13790_ clknet_leaf_83_clk _00903_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08656__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ cpu.f0.write_data\[3\] net499 _01762_ _01768_ vssd1 vssd1 vccd1 vccd1 _01724_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10121__C1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12672_ net2634 cpu.LCD0.row_2\[66\] net1001 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XANTENNA__09409__A2 _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__A _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14411_ clknet_leaf_37_clk _01522_ net1260 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11623_ net2427 net152 net358 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XANTENNA__10694__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__B _05030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__A1 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12475__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_22_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13402__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06744__Y _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14528__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ clknet_leaf_56_clk _01455_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.lcd_rs sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire510 _02793_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_2
XFILLER_0_65_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ net2806 net181 net369 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XANTENNA__10975__A1 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14463__Q cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10505_ net1509 net916 net751 a1.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 _00178_
+ sky130_fd_sc_hd__a22o_1
X_14273_ clknet_leaf_66_clk _01386_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11485_ net2063 net190 net374 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XANTENNA__12177__B1 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09784__A _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ clknet_leaf_89_clk _00404_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ net1125 _01821_ net264 vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__or3_1
XANTENNA__10727__A1 _05016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13552__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07053__C1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ clknet_leaf_53_clk net2403 net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10367_ cpu.f0.i\[28\] net308 _05589_ cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 _05599_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_72_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ net746 _05996_ _05997_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and3_4
X_10298_ cpu.f0.i\[18\] _05534_ _05540_ net307 vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__o211a_1
X_13086_ clknet_leaf_53_clk _00266_ net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_89_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09345__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ cpu.LCD0.cnt_20ms\[13\] cpu.LCD0.cnt_20ms\[12\] cpu.LCD0.cnt_20ms\[11\] cpu.LCD0.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_89_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13988_ clknet_leaf_95_clk _01101_ net1219 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07108__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__B1 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14058__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14638__Q cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12939_ clknet_leaf_28_clk _00128_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08856__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06460_ a1.curr_state\[2\] a1.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__nor2_1
XANTENNA__09959__A cpu.IM0.address_IM\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ clknet_leaf_50_clk net1476 net1382 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09678__B _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06391_ cpu.f0.i\[15\] vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08130_ cpu.RF0.registers\[1\]\[23\] net714 net674 cpu.RF0.registers\[6\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__A0 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08061_ net1087 cpu.RF0.registers\[20\]\[25\] net875 vssd1 vssd1 vccd1 vccd1 _03352_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ cpu.RF0.registers\[10\]\[23\] net569 _02277_ _02287_ _02297_ vssd1 vssd1
+ vccd1 vccd1 _02303_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12168__B1 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap810 _02143_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload38_A clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10194__A2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net934 cpu.RF0.registers\[7\]\[26\] net844 vssd1 vssd1 vccd1 vccd1 _04254_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_51_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08139__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ net958 cpu.RF0.registers\[15\]\[30\] net826 vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10920__X _05834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ cpu.RF0.registers\[10\]\[17\] net691 _04168_ _04170_ _04176_ vssd1 vssd1
+ vccd1 vccd1 _04185_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_32_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1008_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ net1059 cpu.RF0.registers\[31\]\[24\] net828 net598 cpu.RF0.registers\[13\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a32o_1
XANTENNA__07898__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout370_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ cpu.RF0.registers\[8\]\[21\] net611 net588 cpu.RF0.registers\[1\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ net288 _04804_ _04805_ _04802_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_49_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06727_ net1081 cpu.RF0.registers\[28\]\[30\] net867 vssd1 vssd1 vccd1 vccd1 _02018_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ _04086_ net440 _04158_ _04194_ net463 net457 vssd1 vssd1 vccd1 vccd1 _04737_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_45_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06658_ a1.CPU_DAT_O\[26\] net893 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[26\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_26_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08773__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09377_ _03402_ net443 net466 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06589_ cpu.LCD0.cnt_500hz\[7\] cpu.LCD0.cnt_500hz\[6\] cpu.LCD0.cnt_500hz\[9\] cpu.LCD0.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_69_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11403__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08328_ cpu.RF0.registers\[31\]\[12\] net687 _03604_ _03609_ _03611_ vssd1 vssd1
+ vccd1 vccd1 _03619_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_95_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06724__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08259_ cpu.RF0.registers\[28\]\[15\] net706 net648 cpu.RF0.registers\[25\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12159__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ net1677 net237 net400 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__mux2_1
XANTENNA__09024__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ net1471 net729 _05478_ cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__a22o_1
XANTENNA__06740__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__A _02094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _05398_ _05417_ _05416_ _05406_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07050__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10830__X _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ cpu.IM0.address_IM\[20\] _05341_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__nor2_1
Xhold9 net110 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09878__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ clknet_leaf_64_clk _01024_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14200__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09115__Y _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_61_clk _00955_ net1349 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14458__Q cpu.f0.i\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13773_ clknet_leaf_104_clk _00886_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10985_ net273 _05874_ _05875_ net925 a1.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1
+ _00425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08302__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14350__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ net1431 cpu.LCD0.row_2\[118\] net1006 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12655_ net2789 net2691 net1009 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11313__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ net1780 net229 net360 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
X_12586_ net1128 cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ clknet_leaf_56_clk _01438_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ net2669 net248 net369 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09010__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 cpu.RF0.registers\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ clknet_leaf_75_clk _01369_ net1334 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06931__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ net1832 net239 net376 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08369__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ clknet_leaf_93_clk _00387_ net1238 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10419_ net1126 _05627_ net265 net2198 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__a2bb2o_1
X_14187_ clknet_leaf_90_clk _01300_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11399_ net1929 net139 net386 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
X_13138_ clknet_leaf_52_clk net2685 net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11268__B cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11983__S net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13069_ clknet_leaf_52_clk net2517 net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 cpu.RF0.registers\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09869__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13448__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ net964 cpu.RF0.registers\[3\]\[13\] net821 vssd1 vssd1 vccd1 vccd1 _02921_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06378__A cpu.f0.i\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07561_ net1053 cpu.RF0.registers\[21\]\[8\] net797 vssd1 vssd1 vccd1 vccd1 _02852_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09300_ _04370_ _04385_ _04389_ net301 _04382_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o221a_1
X_06512_ cpu.f0.num\[28\] cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07492_ cpu.RF0.registers\[3\]\[5\] net610 _02774_ _02776_ _02778_ vssd1 vssd1 vccd1
+ vccd1 _02783_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_17_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09231_ net464 _04483_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o21a_1
X_06443_ net1118 _01848_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11223__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06374_ cpu.DM0.state\[2\] vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09162_ _03304_ _04293_ _04291_ _03238_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__inv_2
X_09093_ net487 _02681_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__nor2_4
XFILLER_0_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout216_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08044_ cpu.IM0.address_IM\[24\] net553 _03333_ _03334_ vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07280__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold910 cpu.LCD0.row_1\[74\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 a1.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold932 cpu.LCD0.row_2\[59\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold943 cpu.LCD0.row_2\[8\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold954 _01679_ vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold965 _00280_ vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold976 cpu.LCD0.row_2\[112\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13921__RESET_B net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold987 cpu.RF0.registers\[21\]\[29\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 cpu.LCD0.row_2\[104\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net629 _04774_ net931 vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07375__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14223__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_A _02173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ cpu.RF0.registers\[17\]\[27\] net694 net674 cpu.RF0.registers\[6\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__a22o_1
XANTENNA__08768__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07672__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ net1079 cpu.RF0.registers\[16\]\[17\] net841 vssd1 vssd1 vccd1 vccd1 _04168_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08532__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14373__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ _03115_ _03116_ net522 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07740__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ net962 cpu.RF0.registers\[12\]\[21\] net766 vssd1 vssd1 vccd1 vccd1 _03050_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_79_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ net989 cpu.f0.data_adr\[16\] vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08934__C net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09429_ _04669_ _04719_ net455 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11133__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09111__B _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ net2910 net534 vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net1123 net1522 net531 cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 _01497_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ clknet_leaf_83_clk _01223_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ net2860 net172 net394 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
XANTENNA__06751__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A1 _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ clknet_leaf_91_clk _01154_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11253_ net2310 net191 net402 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10158__A2 _05424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ net715 net132 _05466_ net627 vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a31o_1
XANTENNA__13357__Q cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ net2196 net193 net413 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10135_ net625 _05107_ net1022 vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07582__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ net716 net133 _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a21o_1
XANTENNA__09720__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825_ clknet_leaf_67_clk _00938_ net1298 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12607__A1 cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09005__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ clknet_leaf_12_clk _00869_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10968_ _02938_ net515 _05852_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a21o_1
XANTENNA__06926__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ cpu.LCD0.row_2\[109\] cpu.LCD0.row_2\[101\] net998 vssd1 vssd1 vccd1 vccd1
+ _01700_ sky130_fd_sc_hd__mux2_1
XANTENNA__08844__C net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13687_ clknet_leaf_64_clk _00800_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06645__B net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10899_ _05357_ _05818_ net722 vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__mux2_4
XANTENNA__11043__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13890__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ net2285 net2146 net1007 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11978__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ _06333_ net1552 _06320_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09448__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14308_ clknet_leaf_96_clk _01421_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13120__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 a1.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06661__A a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 cpu.RF0.registers\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14246__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold228 _00179_ vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__B1 cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold239 cpu.SR1.char_in\[6\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ clknet_leaf_0_clk _01352_ net1142 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09972__A cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07014__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout708 _02014_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_6
XANTENNA__07195__C net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_2
X_08800_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__inv_2
XANTENNA__11566__X _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12602__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net487 _04762_ _04834_ _04384_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a221o_1
XANTENNA__14396__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ net1027 cpu.RF0.registers\[29\]\[23\] net790 vssd1 vssd1 vccd1 vccd1 _02283_
+ sky130_fd_sc_hd__and3_1
X_08731_ _04010_ _04013_ _04017_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11218__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_2
X_08662_ cpu.RF0.registers\[5\]\[2\] net703 net673 cpu.RF0.registers\[29\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a22o_1
XANTENNA__06525__B2 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ cpu.CU0.funct3\[1\] _02314_ _02313_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__a21o_1
X_08593_ cpu.RF0.registers\[9\]\[4\] net700 net694 cpu.RF0.registers\[17\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a22o_1
X_07544_ net973 cpu.RF0.registers\[10\]\[8\] net788 vssd1 vssd1 vccd1 vccd1 _02835_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__B1 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14191__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06836__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10085__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ net1060 cpu.RF0.registers\[26\]\[5\] net789 vssd1 vssd1 vccd1 vccd1 _02766_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14120__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_A _05938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09214_ net465 net448 _04486_ net453 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__o211a_1
X_06426_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__A1 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11888__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ net462 _03992_ _04026_ net450 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__o211a_1
XANTENNA__08435__D1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06357_ net2420 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__A2 _02543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09076_ _04365_ _04366_ net455 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08027_ net1097 cpu.RF0.registers\[21\]\[24\] net865 vssd1 vssd1 vccd1 vccd1 _03318_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 cpu.LCD0.row_2\[32\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 cpu.RF0.registers\[11\]\[2\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13613__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold762 cpu.RF0.registers\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold773 _00239_ vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__A cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 a1.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 cpu.RF0.registers\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ cpu.IM0.address_IM\[12\] _02869_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__xor2_2
X_08929_ net1084 cpu.RF0.registers\[18\]\[27\] net855 vssd1 vssd1 vccd1 vccd1 _04220_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08929__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13763__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1440 cpu.c0.count\[11\] vssd1 vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 a1.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11940_ net2424 net215 net319 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09106__B _04395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1462 a1.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net2868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 cpu.RF0.registers\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net2879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08010__B _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1484 cpu.RF0.registers\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net2890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1495 cpu.RF0.registers\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net2901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ net1748 net227 net328 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14119__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14208__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ clknet_leaf_100_clk _00723_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10822_ net2368 net558 net536 _05762_ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__a22o_1
X_14590_ clknet_leaf_47_clk _01692_ net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[101\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12100__X _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09122__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ clknet_leaf_9_clk _00654_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10753_ net1613 net559 net537 _05713_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__a22o_1
XANTENNA__10268__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ clknet_leaf_8_clk _00585_ net1161 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13143__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ cpu.LCD0.row_1\[90\] net2311 net897 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XANTENNA__08961__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07492__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14269__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11798__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ net1589 net731 net501 _06235_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__o22a_1
XANTENNA__09776__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12773__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12354_ cpu.K0.enable net1131 cpu.K0.count\[0\] vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07244__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__C_N net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ net2723 net252 net397 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__mux2_1
XANTENNA__13293__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12285_ cpu.LCD0.row_2\[23\] _06003_ _06037_ cpu.LCD0.row_1\[79\] _06178_ vssd1 vssd1
+ vccd1 vccd1 _06179_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ clknet_leaf_99_clk _01137_ net1235 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ net2568 net236 net404 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__mux2_1
XANTENNA__10000__A1 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__B2 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ net2914 net136 net414 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08839__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ cpu.IM0.address_IM\[23\] _05376_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__nor2_1
X_11098_ net2030 net147 net424 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__mux2_1
XANTENNA__11038__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10049_ cpu.IM0.address_IM\[18\] _02349_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10877__S net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__B2 cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13808_ clknet_leaf_74_clk _00921_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06656__A a1.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13739_ clknet_leaf_91_clk _00852_ net1278 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__A cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07260_ net1062 cpu.RF0.registers\[21\]\[7\] net798 vssd1 vssd1 vccd1 vccd1 _02551_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07191_ net970 cpu.RF0.registers\[4\]\[10\] net783 vssd1 vssd1 vccd1 vccd1 _02482_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11501__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13636__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12764__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07918__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14381__Q cpu.IG0.Instr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09901_ cpu.IM0.address_IM\[5\] _05178_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_98_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13786__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload20_A clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _05764_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_2
Xfanout516 _05850_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_4
Xfanout527 _01892_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_2
X_09832_ _03475_ _04552_ _03511_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__a21oi_1
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10542__A2 a1.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_2
X_09763_ _04397_ _04393_ _04999_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__mux2_1
XANTENNA__07653__C _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ net1050 cpu.RF0.registers\[31\]\[25\] net830 net623 vssd1 vssd1 vccd1 vccd1
+ _02266_ sky130_fd_sc_hd__a31o_1
XANTENNA__10360__B cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ cpu.RF0.registers\[14\]\[0\] net649 net643 cpu.RF0.registers\[3\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _04962_ _04984_ _04956_ _04960_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__o211a_1
XANTENNA__09696__B1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08645_ net1102 cpu.RF0.registers\[24\]\[2\] net872 vssd1 vssd1 vccd1 vccd1 _03936_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout548_A _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08576_ net304 _02760_ net492 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08484__C net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14411__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07527_ cpu.RF0.registers\[26\]\[6\] net600 _02175_ cpu.RF0.registers\[6\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09877__A cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06853__X _02144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07458_ cpu.RF0.registers\[26\]\[1\] net599 _02725_ _02731_ _02743_ vssd1 vssd1 vccd1
+ vccd1 _02749_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11007__A0 cpu.f0.write_data\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06409_ cpu.c0.count\[1\] cpu.c0.count\[0\] cpu.c0.count\[3\] cpu.c0.count\[2\] vssd1
+ vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07389_ net524 _02679_ _02645_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11411__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14561__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12755__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ _04417_ _04418_ net456 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__mux2_1
XANTENNA__09620__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08974__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ cpu.RF0.registers\[1\]\[31\] net588 _04333_ _04335_ _04343_ vssd1 vssd1 vccd1
+ vccd1 _04350_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12070_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 cpu.RF0.registers\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 cpu.RF0.registers\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 cpu.f0.data_adr\[18\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _03192_ net533 net283 vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08726__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08021__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ clknet_leaf_28_clk net1519 net1183 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09687__B1 _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A2 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 cpu.RF0.registers\[0\]\[26\] vssd1 vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13509__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11923_ net2896 net157 net322 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
Xhold1281 cpu.RF0.registers\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 cpu.RF0.registers\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
X_14642_ clknet_leaf_23_clk _01743_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11854_ net2859 net152 net330 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14091__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14466__Q cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ cpu.IM0.address_IM\[26\] net1013 net284 _05750_ vssd1 vssd1 vccd1 vccd1 _05751_
+ sky130_fd_sc_hd__a22o_1
X_14573_ clknet_leaf_49_clk _01675_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[84\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ net2320 net181 net341 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13524_ clknet_leaf_69_clk _00637_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10736_ net1602 net559 net537 _05701_ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__a22o_1
XANTENNA__07465__A2 _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__X _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13455_ clknet_leaf_80_clk _00568_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ net2737 net2607 net906 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11321__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ cpu.DM0.readdata\[11\] net732 _06226_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13386_ clknet_leaf_102_clk _00499_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ cpu.LCD0.row_1\[4\] cpu.LCD0.row_1\[12\] net899 vssd1 vssd1 vccd1 vccd1 _00228_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__10221__B2 cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12337_ _06208_ _06209_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__nor2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__10772__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ cpu.LCD0.row_1\[62\] _06025_ _06028_ cpu.LCD0.row_1\[118\] _06162_ vssd1
+ vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09953__C cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13039__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A1 _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ clknet_leaf_64_clk _01120_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11219_ net1944 net207 net406 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
X_12199_ cpu.LCD0.row_1\[3\] _06015_ _06019_ cpu.LCD0.row_1\[51\] _06096_ vssd1 vssd1
+ vccd1 vccd1 _06097_ sky130_fd_sc_hd__a221o_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__07386__D1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07473__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06760_ net948 net842 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__nand2_4
XANTENNA__14434__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06691_ net1594 net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[27\] sky130_fd_sc_hd__and2_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ cpu.RF0.registers\[11\]\[9\] net690 net674 cpu.RF0.registers\[6\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06386__A cpu.f0.i\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08361_ cpu.RF0.registers\[13\]\[11\] net659 net650 cpu.RF0.registers\[14\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14584__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ net523 _02583_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__nand2_2
XFILLER_0_74_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09697__A _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07456__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ cpu.RF0.registers\[12\]\[13\] net696 net677 cpu.RF0.registers\[4\]\[13\]
+ _03570_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07243_ cpu.RF0.registers\[3\]\[9\] net609 _02516_ _02521_ _02524_ vssd1 vssd1 vccd1
+ vccd1 _02534_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12737__A0 cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07208__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ _02461_ _02462_ _02463_ _02464_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_41_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09602__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__A2 _05986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10923__X _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09905__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08708__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 _05943_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_4
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_8
Xfanout335 _05937_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11712__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 net349 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_6
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _04414_ _04860_ _05105_ _04480_ _05104_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a221o_1
Xfanout357 _05932_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout368 _05929_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_8
Xfanout379 net381 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_6
XANTENNA_fanout665_A _02050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09746_ net458 _04908_ _05036_ _02758_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__o211a_1
XANTENNA__12268__A2 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06958_ net525 _02247_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__or2_1
XANTENNA__06848__X _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09224__X _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09677_ net306 _03899_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nor2_1
X_06889_ net1038 cpu.RF0.registers\[18\]\[27\] net770 vssd1 vssd1 vccd1 vccd1 _02180_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout832_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ cpu.RF0.registers\[5\]\[3\] net704 net698 cpu.RF0.registers\[12\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13801__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06727__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12448__D net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net1105 cpu.RF0.registers\[26\]\[5\] _02025_ vssd1 vssd1 vccd1 vccd1 _03850_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ net1967 net245 net365 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ net67 net919 vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__and2_1
XANTENNA__13951__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13435__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12728__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ clknet_leaf_37_clk _00420_ net1258 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10452_ net32 net755 _05640_ a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08016__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08947__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11929__X _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ clknet_leaf_37_clk _00351_ net1264 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10383_ net1124 _05609_ net266 net2140 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10833__X _05772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14307__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12122_ cpu.LCD0.row_1\[88\] _06021_ _06022_ cpu.LCD0.row_2\[120\] vssd1 vssd1 vccd1
+ vccd1 _06023_ sky130_fd_sc_hd__a22o_1
XANTENNA__07855__A _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07080__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08303__X _03594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ cpu.LCD0.cnt_500hz\[5\] _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14294__RESET_B net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ cpu.f0.write_data\[23\] _05888_ net985 vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14457__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout880 _02008_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_8
Xfanout891 _01951_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_2
XANTENNA__12259__A2 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ clknet_leaf_20_clk _00144_ net1169 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11316__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ net2268 net217 net322 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12886_ clknet_leaf_29_clk _00007_ net1201 vssd1 vssd1 vccd1 vccd1 cpu.f0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_73_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07686__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14625_ clknet_leaf_30_clk _01726_ net1203 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10690__A1 cpu.LCD0.row_1\[104\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ net1902 net231 net333 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__mux2_1
XANTENNA__09013__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ clknet_leaf_46_clk _01658_ net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11768_ net2071 net247 net340 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__mux2_1
XANTENNA__06934__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08852__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ net993 _05058_ net285 net1014 cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1
+ _05690_ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13507_ clknet_leaf_74_clk _00620_ net1317 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14487_ clknet_leaf_57_clk _01590_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11699_ net1618 net239 net348 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11051__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap1131 _01996_ vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_2
X_13438_ clknet_leaf_85_clk _00551_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11986__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10890__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13369_ clknet_leaf_42_clk _00482_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10745__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ cpu.RF0.registers\[1\]\[30\] net588 net576 cpu.RF0.registers\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a22o_1
XANTENNA__10191__A cpu.IM0.address_IM\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ cpu.RF0.registers\[9\]\[28\] net574 net565 cpu.RF0.registers\[30\]\[28\]
+ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10902__C1 _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ _02830_ _03833_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
XANTENNA__08571__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06812_ net1118 _01846_ _02083_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13824__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07792_ net1031 cpu.RF0.registers\[23\]\[22\] net816 vssd1 vssd1 vccd1 vccd1 _03083_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09531_ _03664_ _03698_ net468 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06743_ net936 cpu.RF0.registers\[15\]\[30\] net859 vssd1 vssd1 vccd1 vccd1 _02034_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06828__B _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ net493 _04664_ _04735_ _04743_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a311oi_4
X_06674_ a1.CPU_DAT_O\[10\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[10\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ net1079 cpu.RF0.registers\[20\]\[9\] net874 vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13974__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _04617_ _04639_ _04663_ _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_47_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout246_A _05776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ _03540_ _03568_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07429__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08275_ _02436_ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout413_A _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13204__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07226_ net1034 cpu.RF0.registers\[21\]\[9\] net795 vssd1 vssd1 vccd1 vccd1 _02517_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07157_ net1043 cpu.RF0.registers\[25\]\[11\] net757 vssd1 vssd1 vccd1 vccd1 _02448_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_93_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1322_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13354__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07601__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ cpu.RF0.registers\[8\]\[18\] net612 _02378_ net622 vssd1 vssd1 vccd1 vccd1
+ _02379_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout782_A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1430_A cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12489__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_2
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
Xfanout143 _05841_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 _05827_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
Xfanout176 _05807_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout198 net200 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09729_ _04429_ _04438_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12740_ cpu.f0.i\[3\] _01871_ _06332_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12671_ net2471 cpu.LCD0.row_2\[65\] net1009 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14410_ clknet_leaf_35_clk net1630 net1252 vssd1 vssd1 vccd1 vccd1 cpu.DM0.readdata\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11622_ net2871 net163 net358 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06754__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__C _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_52_clk _01454_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11553_ net1570 net170 net366 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08093__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__A2 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10504_ net1438 net918 net750 a1.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 _00177_
+ sky130_fd_sc_hd__a22o_1
X_14272_ clknet_leaf_3_clk _01385_ net1160 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07840__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ cpu.RF0.registers\[14\]\[16\] net206 net374 vssd1 vssd1 vccd1 vccd1 _00904_
+ sky130_fd_sc_hd__mux2_1
X_13223_ clknet_leaf_100_clk _00403_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ _01819_ net270 _05635_ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09784__B _04881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06760__Y _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07585__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ clknet_leaf_52_clk _00334_ net1372 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10366_ net1537 net726 _05598_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ net745 _05984_ _05989_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and3_4
X_13085_ clknet_leaf_51_clk net2366 net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ cpu.f0.i\[18\] _05534_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__nand2_1
XANTENNA__13847__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__C net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12036_ cpu.LCD0.cnt_20ms\[9\] cpu.LCD0.cnt_20ms\[7\] cpu.LCD0.cnt_20ms\[6\] cpu.LCD0.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__or4b_1
XFILLER_0_40_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09008__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06929__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08847__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13997__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ clknet_leaf_79_clk _01100_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11046__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ clknet_leaf_28_clk _00127_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_76_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10738__X _05703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09959__B cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ clknet_leaf_5_clk cpu.c0.next_count\[0\] net1145 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13227__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14608_ clknet_leaf_52_clk net2440 net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08608__A1 cpu.IM0.address_IM\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06390_ cpu.f0.num\[15\] vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06664__A a1.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09805__B1 _05095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14539_ clknet_leaf_61_clk _01641_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08060_ net943 cpu.RF0.registers\[13\]\[25\] net850 vssd1 vssd1 vccd1 vccd1 _03351_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13377__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07198__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14622__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07011_ cpu.RF0.registers\[7\]\[23\] net596 _02289_ _02294_ _02295_ vssd1 vssd1 vccd1
+ vccd1 _02302_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12605__S net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__B1 cpu.IM0.address_IM\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07044__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07926__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14145__RESET_B net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ net1080 cpu.RF0.registers\[27\]\[26\] net880 vssd1 vssd1 vccd1 vccd1 _04253_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07913_ net1029 cpu.RF0.registers\[26\]\[30\] net787 vssd1 vssd1 vccd1 vccd1 _03204_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ cpu.RF0.registers\[8\]\[17\] net708 _04169_ _04172_ _04174_ vssd1 vssd1 vccd1
+ vccd1 _04184_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_32_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout196_A _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _03128_ _03130_ _03132_ _03134_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14002__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07661__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ cpu.RF0.registers\[19\]\[21\] net616 _03058_ _03063_ _03064_ vssd1 vssd1
+ vccd1 vccd1 _03066_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout363_A _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ net296 net293 _04803_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__mux2_1
X_06726_ net1092 net868 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ _04158_ _04194_ net463 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06657_ net1858 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[25\] sky130_fd_sc_hd__and2_1
XANTENNA_fanout530_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14152__CLK clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09376_ _04089_ _04665_ _04127_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__o21ai_1
X_06588_ cpu.LCD0.cnt_500hz\[5\] cpu.LCD0.cnt_500hz\[8\] cpu.LCD0.cnt_500hz\[11\]
+ cpu.LCD0.cnt_500hz\[4\] vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_23_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07022__X _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08327_ cpu.RF0.registers\[18\]\[12\] net680 net653 cpu.RF0.registers\[7\]\[12\]
+ _03603_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09272__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A2 _02037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08258_ cpu.RF0.registers\[11\]\[15\] net688 net671 cpu.RF0.registers\[23\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07822__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12159__A1 cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07209_ cpu.RF0.registers\[7\]\[10\] net595 _02486_ _02490_ _02494_ vssd1 vssd1 vccd1
+ vccd1 _02500_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08189_ net1088 cpu.RF0.registers\[19\]\[21\] net835 vssd1 vssd1 vccd1 vccd1 _03480_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10824__A cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ cpu.f0.data_adr\[4\] net729 _05478_ cpu.f0.i\[2\] vssd1 vssd1 vccd1 vccd1
+ _00057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10543__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__Q cpu.IM0.address_IM\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _05398_ _05417_ _05406_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__o21a_1
XANTENNA__10590__A0 _05683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ cpu.IM0.address_IM\[20\] _05341_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08535__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ clknet_leaf_57_clk _01023_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12103__X _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__B1 cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ clknet_leaf_76_clk _00954_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13772_ clknet_leaf_88_clk _00885_ net1295 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net985 cpu.f0.write_data\[17\] vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12723_ cpu.LCD0.row_2\[125\] cpu.LCD0.row_2\[117\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12654_ net2186 cpu.LCD0.row_2\[48\] net1010 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__mux2_1
XANTENNA__06484__A cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12398__A1 cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14474__Q cpu.SR1.char_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14645__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11605_ net1834 net234 net360 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
X_12585_ _06346_ net1645 _06320_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux2_1
XANTENNA__08066__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ net2815 net252 net369 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
X_14324_ clknet_leaf_57_clk _01437_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06771__X _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14255_ clknet_leaf_82_clk _01368_ net1285 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ _05766_ net503 _05912_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__and3_4
XFILLER_0_81_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13206_ clknet_leaf_91_clk _00386_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ cpu.f0.i\[21\] net269 vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__nand2_1
X_14186_ clknet_leaf_100_clk _01299_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11398_ cpu.RF0.registers\[11\]\[29\] net143 net388 vssd1 vssd1 vccd1 vccd1 _00821_
+ sky130_fd_sc_hd__mux2_1
X_13137_ clknet_leaf_48_clk _00317_ net1355 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10349_ _05582_ _05583_ net526 vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10581__A0 cpu.f0.write_data\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ clknet_leaf_49_clk _00248_ net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10381__A1_N net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14025__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09869__A3 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ net2894 net152 net310 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10333__B1 _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14649__Q cpu.f0.write_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07481__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ cpu.RF0.registers\[23\]\[8\] net613 net607 cpu.RF0.registers\[24\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06511_ cpu.f0.num\[13\] cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_0_clk_X clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07491_ cpu.RF0.registers\[6\]\[5\] net583 net567 cpu.RF0.registers\[11\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11504__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ net453 _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nand2_1
X_06442_ cpu.CU0.opcode\[4\] _01847_ net1118 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__nor3b_2
XANTENNA__06515__A2_N net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06394__A cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14384__Q cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _01781_ _04450_ _04448_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__mux2_1
XANTENNA__12389__B2 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06373_ net1 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10939__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08112_ _03118_ _03122_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09092_ net305 _04381_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload50_A clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ cpu.RF0.registers\[0\]\[24\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__o21a_1
Xhold900 cpu.LCD0.row_2\[99\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 _00298_ vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06841__B net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold922 cpu.RF0.registers\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold933 _01650_ vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08114__A _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold944 cpu.RF0.registers\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold955 cpu.RF0.registers\[28\]\[17\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 cpu.RF0.registers\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _01703_ vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold988 cpu.LCD0.row_2\[97\] vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net126 _05273_ _05270_ net629 vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a211o_1
Xhold999 _01695_ vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07953__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _04232_ _04233_ _04234_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout578_A _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ net1076 cpu.RF0.registers\[27\]\[17\] net880 vssd1 vssd1 vccd1 vccd1 _04167_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10324__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10875__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ net546 _03116_ _03117_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_93_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07758_ net1042 cpu.RF0.registers\[23\]\[21\] net817 vssd1 vssd1 vccd1 vccd1 _03049_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06709_ cpu.CU0.opcode\[1\] cpu.CU0.opcode\[0\] cpu.CU0.opcode\[2\] vssd1 vssd1 vccd1
+ vccd1 _02000_ sky130_fd_sc_hd__and3_1
XANTENNA__13542__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout912_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _02971_ _02977_ _02978_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__or4_1
XANTENNA__08296__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1275_X net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09428_ net441 net439 net467 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12807__Q cpu.IM0.address_IM\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ net452 _04372_ _04387_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a31o_2
XANTENNA__13692__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ net1123 net1593 net531 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 _01496_
+ sky130_fd_sc_hd__a22o_1
X_11321_ net2840 net187 net396 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06751__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ clknet_leaf_19_clk _01153_ net1180 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09548__A2 _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net2741 _05810_ net402 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08024__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__A1 cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _05464_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ net1687 net199 net410 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__mux2_1
XANTENNA__08959__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__X _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ net125 _05400_ _05402_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08508__B1 _02122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13072__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06782__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _05337_ _05338_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__xor2_1
XANTENNA__06479__A cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10315__B1 cpu.f0.i\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13824_ clknet_leaf_5_clk _00937_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10967_ net276 _05861_ _05862_ net928 net2085 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a32o_1
X_13755_ clknet_leaf_12_clk _00868_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11324__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ cpu.LCD0.row_2\[108\] cpu.LCD0.row_2\[100\] net1008 vssd1 vssd1 vccd1 vccd1
+ _01699_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13686_ clknet_leaf_59_clk _00799_ net1348 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10898_ cpu.DM0.readdata\[20\] _05096_ net738 vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ net2448 net2588 net1007 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
XANTENNA__08039__A2 _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12240__B1 _06033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ net1128 cpu.DM0.data_i\[3\] _06307_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06942__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14307_ clknet_leaf_79_clk _01420_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11519_ net2334 net188 net371 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__mux2_1
X_12499_ _05527_ _06268_ _06282_ cpu.f0.i\[16\] net262 vssd1 vssd1 vccd1 vccd1 _01564_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 a1.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06661__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold218 cpu.LCD0.row_1\[121\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 cpu.RF0.registers\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ clknet_leaf_84_clk _01351_ net1270 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07476__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13415__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ clknet_leaf_91_clk _01282_ net1240 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08211__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08869__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_6
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07773__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ net1027 cpu.RF0.registers\[24\]\[23\] net811 vssd1 vssd1 vccd1 vccd1 _02282_
+ sky130_fd_sc_hd__and3_1
X_08730_ cpu.RF0.registers\[7\]\[0\] net652 _04018_ _04019_ _04020_ vssd1 vssd1 vccd1
+ vccd1 _04021_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06389__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1280 net1283 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__clkbuf_2
X_08661_ cpu.RF0.registers\[9\]\[2\] net701 net637 cpu.RF0.registers\[16\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a22o_1
Xfanout1291 net1300 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_2
XANTENNA__13565__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07612_ net522 _02901_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__o21ai_4
X_08592_ net948 cpu.RF0.registers\[15\]\[4\] net857 vssd1 vssd1 vccd1 vccd1 _03883_
+ sky130_fd_sc_hd__and3_1
X_07543_ net973 cpu.RF0.registers\[1\]\[8\] net806 vssd1 vssd1 vccd1 vccd1 _02834_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08278__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06836__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_A _05832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11234__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ net1056 cpu.RF0.registers\[30\]\[5\] net764 vssd1 vssd1 vccd1 vccd1 _02765_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _04500_ _04503_ net470 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__mux2_1
X_06425_ cpu.c0.count\[9\] _01835_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout326_A _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net462 _03992_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__nor2_1
XANTENNA__12231__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06356_ cpu.LCD0.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ net441 net440 net466 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1235_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ net1097 cpu.RF0.registers\[30\]\[24\] net840 vssd1 vssd1 vccd1 vccd1 _03317_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold730 cpu.RF0.registers\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _01623_ vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout695_A _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13095__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 cpu.RF0.registers\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__B _02583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold763 cpu.RF0.registers\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 cpu.RF0.registers\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 cpu.RF0.registers\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 cpu.RF0.registers\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08779__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ cpu.IM0.address_IM\[11\] _05258_ net1023 vssd1 vssd1 vccd1 vccd1 _00034_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13908__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10560__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net1083 cpu.RF0.registers\[20\]\[27\] net874 vssd1 vssd1 vccd1 vccd1 _04219_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09163__A0 _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1430 cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10848__A1 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1441 cpu.RF0.registers\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1452 cpu.c0.count\[12\] vssd1 vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14490__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ _04146_ _04147_ _04148_ _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__or4_1
Xhold1463 cpu.RF0.registers\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1474 cpu.RF0.registers\[30\]\[6\] vssd1 vssd1 vccd1 vccd1 net2880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 cpu.RF0.registers\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net2891 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12932__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1496 cpu.RF0.registers\[0\]\[2\] vssd1 vssd1 vccd1 vccd1 net2902 sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ net2776 net228 net328 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06586__X _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ cpu.IM0.address_IM\[31\] net1013 net284 _05761_ vssd1 vssd1 vccd1 vccd1 _05762_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06746__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ cpu.IM0.address_IM\[11\] net1015 net286 _05712_ vssd1 vssd1 vccd1 vccd1 _05713_
+ sky130_fd_sc_hd__a22o_1
X_13540_ clknet_leaf_96_clk _00653_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08019__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14248__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ clknet_leaf_106_clk _00584_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ net2508 cpu.LCD0.row_1\[97\] net911 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
XANTENNA__10836__X _05774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11025__A1 _05902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12422_ cpu.DM0.data_i\[19\] net535 vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__and2_1
XANTENNA__12222__B1 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06762__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ cpu.K0.enable cpu.K0.count\[0\] net1131 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__and3_1
XANTENNA__10784__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ net2784 net254 net397 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__mux2_1
X_12284_ cpu.LCD0.row_1\[7\] _06015_ _06034_ cpu.LCD0.row_2\[31\] vssd1 vssd1 vccd1
+ vccd1 _06178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12525__A1 cpu.f0.i\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ clknet_leaf_82_clk _01136_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09926__C1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ _05765_ net504 _05915_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__and3_4
XANTENNA__12703__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net2225 net142 net415 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__mux2_1
XANTENNA__11319__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ cpu.IM0.address_IM\[23\] _05376_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__and2_2
XANTENNA__12289__B1 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ net1851 net150 net422 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
X_10048_ cpu.IM0.address_IM\[17\] net930 _05322_ _05323_ vssd1 vssd1 vccd1 vccd1 _00040_
+ sky130_fd_sc_hd__a22o_1
Xhold90 net80 vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06937__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__A2 cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ clknet_leaf_83_clk _00920_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09457__B2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11054__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11999_ net1716 net246 net313 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ clknet_leaf_95_clk _00851_ net1218 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__B cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14213__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10893__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ clknet_leaf_103_clk _00782_ net1158 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09459__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07190_ net1051 cpu.RF0.registers\[29\]\[10\] net793 vssd1 vssd1 vccd1 vccd1 _02481_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06672__A a1.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08590__C _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12764__B2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14363__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _05186_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10922__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout506 _05764_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__dlymetal6s2s_1
X_09831_ _03475_ _03511_ _04552_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and3_1
Xfanout528 _01892_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_2
Xfanout539 _05687_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_2
XANTENNA_clkload13_A clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11229__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ _03995_ _03996_ _04026_ net513 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a31o_1
X_06974_ cpu.RF0.registers\[3\]\[25\] net609 net583 cpu.RF0.registers\[6\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
XANTENNA__12955__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07653__D _02940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08713_ cpu.RF0.registers\[13\]\[0\] net657 net655 cpu.RF0.registers\[2\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a22o_1
X_09693_ _04971_ _04979_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08499__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09696__A1 _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout276_A _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net1102 cpu.RF0.registers\[22\]\[2\] _02038_ vssd1 vssd1 vccd1 vccd1 _03935_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06847__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ cpu.IM0.address_IM\[5\] net554 _03864_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_
+ sky130_fd_sc_hd__a22o_2
XANTENNA__10369__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_A _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07526_ net1058 cpu.RF0.registers\[31\]\[6\] net828 vssd1 vssd1 vccd1 vccd1 _02817_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_77_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11899__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07457_ _02744_ _02745_ _02746_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__or4_1
XANTENNA__09877__B cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1352_A net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06408_ net1927 _01822_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[2\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07388_ cpu.RF0.registers\[0\]\[2\] net619 _02676_ _02678_ vssd1 vssd1 vccd1 vccd1
+ _02679_ sky130_fd_sc_hd__o22a_4
X_09127_ _03534_ net300 net467 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XANTENNA__12755__B2 cpu.f0.i\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10230__A2 cpu.f0.i\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ cpu.RF0.registers\[7\]\[31\] net596 _04325_ _04328_ _04339_ vssd1 vssd1 vccd1
+ vccd1 _04349_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_62_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13730__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _03298_ _03299_ cpu.IM0.address_IM\[28\] net554 vssd1 vssd1 vccd1 vccd1 _03300_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10781__A3 _05733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 cpu.FetchedInstr\[0\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 a1.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A0 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ net2033 net928 net276 _05899_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold582 cpu.RF0.registers\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 cpu.f0.num\[16\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11139__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__Q cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13880__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ clknet_leaf_44_clk net1470 net1304 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
Xhold1260 cpu.RF0.registers\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1271 cpu.FetchedInstr\[7\] vssd1 vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09404__Y _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net2821 net159 net322 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
Xhold1282 cpu.RF0.registers\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12111__X _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1293 cpu.RF0.registers\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06757__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13110__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14236__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14641_ clknet_leaf_23_clk _01742_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_11853_ net1611 net166 net331 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
XANTENNA__09439__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ cpu.f0.data_adr\[26\] _04640_ net989 vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__mux2_1
X_14572_ clknet_leaf_46_clk net1756 net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_11784_ net2094 net170 net338 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__A1 cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13523_ clknet_leaf_69_clk _00636_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ cpu.IM0.address_IM\[6\] net1015 net286 _05700_ vssd1 vssd1 vccd1 vccd1 _05701_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13260__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__A cpu.f0.i\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14386__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11602__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14011__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07588__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ net2805 net2720 net910 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
X_13454_ clknet_leaf_1_clk _00567_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07870__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12828__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06923__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12405_ cpu.DM0.data_i\[11\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13385_ clknet_leaf_103_clk _00498_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ cpu.LCD0.row_1\[3\] net2295 net900 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09611__B2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_49_1697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12336_ net2716 _06207_ net1368 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06976__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12267_ cpu.LCD0.row_2\[6\] _06016_ _06021_ cpu.LCD0.row_1\[94\] vssd1 vssd1 vccd1
+ vccd1 _06162_ sky130_fd_sc_hd__a22o_1
XANTENNA__12978__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10509__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ net2078 net176 net408 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
X_14006_ clknet_leaf_58_clk _01119_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12198_ cpu.LCD0.row_2\[83\] _05990_ _06003_ cpu.LCD0.row_2\[19\] vssd1 vssd1 vccd1
+ vccd1 _06096_ sky130_fd_sc_hd__a22o_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11049__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__10524__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ net2901 net210 net417 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XANTENNA__09127__A0 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08335__D1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ a1.CPU_DAT_O\[26\] net888 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[26\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06667__A a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08585__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09978__A cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13603__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ _03648_ _03649_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08882__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ cpu.RF0.registers\[0\]\[4\] net618 _02598_ _02601_ vssd1 vssd1 vccd1 vccd1
+ _02602_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ cpu.RF0.registers\[14\]\[13\] net650 _03579_ _03580_ _03581_ vssd1 vssd1
+ vccd1 vccd1 _03582_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09697__B _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10476__X _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11512__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ cpu.RF0.registers\[30\]\[9\] net565 _02511_ _02514_ _02532_ vssd1 vssd1 vccd1
+ vccd1 _02533_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07861__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12737__A1 _06329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13753__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ cpu.RF0.registers\[10\]\[11\] net569 _02442_ _02444_ _02446_ vssd1 vssd1
+ vccd1 vccd1 _02464_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_41_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07613__B1 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13734__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06967__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14109__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 _05942_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_6
XANTENNA__07664__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout325 _05940_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout336 _05937_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_6
X_09814_ _04482_ _04853_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__nand2_1
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_8
Xfanout358 _05931_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_8
XANTENNA_fanout1100_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__A0 _05424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _05929_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_4
XANTENNA__13133__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14259__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ net458 _04906_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ cpu.IG0.Instr\[26\] net634 _02210_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout658_A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ _02794_ _03866_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__xor2_2
X_06888_ net1049 net771 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__and2_1
XANTENNA__12298__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ _03915_ _03916_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or3_1
XANTENNA__10099__A cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13283__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06864__X _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ net1105 cpu.RF0.registers\[23\]\[5\] net846 vssd1 vssd1 vccd1 vccd1 _03849_
+ sky130_fd_sc_hd__and3_1
X_07509_ net1057 cpu.RF0.registers\[27\]\[6\] net778 vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10987__A0 cpu.f0.write_data\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ net1107 cpu.RF0.registers\[31\]\[7\] net858 vssd1 vssd1 vccd1 vccd1 _03780_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11422__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ net1134 net2842 net914 _05647_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07852__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__Q cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06743__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07201__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ net31 net753 net563 net2672 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__o22a_1
XANTENNA__10739__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13170_ clknet_leaf_36_clk _00350_ net1263 vssd1 vssd1 vccd1 vccd1 a1.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10382_ cpu.f0.i\[3\] net270 vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ net746 _05987_ net557 vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__and3_4
XANTENNA__12106__X _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net502 _05962_ _05963_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__and3_1
Xhold390 cpu.RF0.registers\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10281__B cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11003_ _02309_ net532 net282 vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_70_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08967__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net873 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
Xfanout881 _02008_ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06758__Y _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13626__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_20_clk _00143_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07135__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 cpu.RF0.registers\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ net2692 net220 net324 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
X_12885_ clknet_leaf_1_clk cpu.c0.next_count\[16\] net1139 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14624_ clknet_leaf_29_clk _01725_ net1203 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06774__X _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net1955 net234 net333 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13776__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08096__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ clknet_leaf_61_clk _01657_ net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10737__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net1669 net251 net341 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__mux2_1
XANTENNA__08635__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13506_ clknet_leaf_10_clk _00619_ net1221 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ net1617 net560 net538 _05689_ vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14486_ clknet_leaf_41_clk _01589_ net1267 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ net505 _05910_ _05915_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13437_ clknet_leaf_89_clk _00550_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ net2333 net2111 net902 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12195__A2 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13368_ clknet_leaf_18_clk _00481_ net1192 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06949__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12319_ net1369 _05949_ _06198_ _05957_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a31o_1
X_13299_ clknet_leaf_34_clk cpu.RU0.next_FetchedData\[6\] net1248 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13156__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09038__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07484__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10191__B _05443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ cpu.RF0.registers\[20\]\[28\] net594 net589 cpu.RF0.registers\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_79_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08877__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__B1 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ cpu.CU0.opcode\[3\] _02091_ net629 net741 net633 vssd1 vssd1 vccd1 vccd1
+ _02102_ sky130_fd_sc_hd__a2111o_2
X_07791_ net957 cpu.RF0.registers\[12\]\[22\] net765 vssd1 vssd1 vccd1 vccd1 _03082_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11507__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09530_ _04603_ _04820_ net470 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__mux2_1
X_06742_ net940 net859 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_30_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06397__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09461_ _04677_ _04710_ _04749_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o211ai_2
XANTENNA__14387__Q cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06673_ a1.CPU_DAT_O\[9\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_94_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08412_ cpu.RF0.registers\[28\]\[9\] net705 net672 cpu.RF0.registers\[29\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__a22o_1
X_09392_ net493 _04666_ _04667_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_47_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08343_ _03601_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout141_A _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09823__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06844__B net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11242__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08274_ net490 _02410_ _03536_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__o21a_1
XANTENNA__07834__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13915__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07659__C net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08117__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07225_ net1034 cpu.RF0.registers\[18\]\[9\] net769 vssd1 vssd1 vccd1 vccd1 _02516_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07021__A _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09587__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07956__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ net1050 cpu.RF0.registers\[27\]\[11\] net777 vssd1 vssd1 vccd1 vccd1 _02447_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06860__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10382__A cpu.f0.i\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07087_ cpu.RF0.registers\[23\]\[18\] net613 net565 cpu.RF0.registers\[30\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1315_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07394__C net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14081__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 cpu.IG0.Instr\[19\] vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout133 net135 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
XANTENNA__13649__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout144 _05839_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XANTENNA__06859__X _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout155 net158 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout166 _05825_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
Xfanout177 net180 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
Xfanout188 _05814_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout942_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ net1092 cpu.RF0.registers\[22\]\[28\] net852 vssd1 vssd1 vccd1 vccd1 _03280_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11417__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _04428_ _04432_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07117__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13799__CLK clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _04802_ _04803_ _04946_ _04948_ _04768_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__o2111ai_2
XANTENNA__10121__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ net2352 net2280 net1009 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09411__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ net2570 net167 net359 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
XANTENNA__13029__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__D _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06754__B net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ clknet_leaf_56_clk _01453_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09130__B _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ net2258 net185 net368 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
XANTENNA__07825__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08027__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ net89 net922 net747 net1481 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__a22o_1
X_11483_ net2139 net174 net376 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
X_14271_ clknet_leaf_106_clk _01384_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13179__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ net266 net1124 cpu.f0.i\[29\] vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__or3b_1
X_13222_ clknet_leaf_103_clk _00402_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06770__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13153_ clknet_leaf_48_clk _00333_ net1355 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[117\]
+ sky130_fd_sc_hd__dfstp_1
X_10365_ net527 _05593_ _05594_ _05597_ net728 vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a311o_1
XANTENNA__08250__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ cpu.LCD0.row_2\[16\] _06003_ _06004_ cpu.LCD0.row_2\[32\] vssd1 vssd1 vccd1
+ vccd1 _06005_ sky130_fd_sc_hd__a22o_1
X_13084_ clknet_leaf_50_clk _00264_ net1382 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ cpu.f0.i\[17\] cpu.f0.i\[18\] _05526_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and3_1
X_12035_ net1660 _05948_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nand2_1
XANTENNA__14574__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11327__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13986_ clknet_leaf_11_clk _01099_ net1224 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08984__X _04275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__A1 _02832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__A2 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ clknet_leaf_29_clk _00126_ net1202 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08856__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06945__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12868_ clknet_leaf_5_clk cpu.c0.next_atmax net1145 vssd1 vssd1 vccd1 vccd1 cpu.K0.enable
+ sky130_fd_sc_hd__dfrtp_1
X_14607_ clknet_leaf_55_clk net2239 net1367 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_11819_ net1854 net168 net335 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
XANTENNA__09805__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06664__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11062__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ cpu.RF0.registers\[0\]\[25\] vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13397__RESET_B net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14538_ clknet_leaf_51_clk _01640_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07479__C net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__A1 cpu.IG0.Instr\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469_ clknet_leaf_22_clk _01579_ net1172 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07292__B2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07010_ cpu.RF0.registers\[12\]\[23\] net572 _02282_ _02283_ _02284_ vssd1 vssd1
+ vccd1 vccd1 _02301_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12168__A2 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__A1 cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap834 _02126_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09991__A cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08961_ net1077 cpu.RF0.registers\[21\]\[26\] net866 vssd1 vssd1 vccd1 vccd1 _04252_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07912_ net1030 cpu.RF0.registers\[28\]\[30\] net765 vssd1 vssd1 vccd1 vccd1 _03203_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12621__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08892_ cpu.RF0.registers\[1\]\[17\] net714 net638 cpu.RF0.registers\[26\]\[17\]
+ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__a221o_1
XANTENNA__07347__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07843_ cpu.RF0.registers\[19\]\[24\] net615 net581 cpu.RF0.registers\[16\]\[24\]
+ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a221o_1
XANTENNA__07898__A3 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13941__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__RESET_B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ net967 cpu.RF0.registers\[5\]\[21\] net796 vssd1 vssd1 vccd1 vccd1 _03065_
+ sky130_fd_sc_hd__and3_1
X_09513_ _02903_ net435 vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06725_ net1114 net1116 net1110 net1112 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_49_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _04055_ _04056_ _04165_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_45_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06656_ a1.CPU_DAT_O\[24\] net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06855__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08773__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ _04089_ _04127_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__or3_1
X_06587_ cpu.LCD0.cnt_500hz\[13\] cpu.LCD0.cnt_500hz\[12\] cpu.LCD0.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout523_A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1265_A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08326_ _03605_ _03614_ _03615_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_95_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14447__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08257_ cpu.RF0.registers\[3\]\[15\] net643 net667 vssd1 vssd1 vccd1 vccd1 _03548_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11700__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12159__A2 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07208_ cpu.RF0.registers\[30\]\[10\] net565 _02482_ _02483_ _02485_ vssd1 vssd1
+ vccd1 vccd1 _02499_ sky130_fd_sc_hd__a2111o_1
X_08188_ net1084 cpu.RF0.registers\[21\]\[21\] net866 vssd1 vssd1 vccd1 vccd1 _03479_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09024__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__B _05763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ cpu.RF0.registers\[3\]\[15\] net609 net599 cpu.RF0.registers\[26\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a22o_1
XANTENNA__08232__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13471__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14597__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11001__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ cpu.IM0.address_IM\[25\] _02272_ _03143_ cpu.IM0.address_IM\[24\] vssd1 vssd1
+ vccd1 vccd1 _05417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10590__A1 cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ net716 net133 _05352_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_7_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08310__A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__A1 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_75_clk _00953_ net1336 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09125__B _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13771_ clknet_leaf_89_clk _00884_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10839__X _05776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ net282 _05873_ net986 vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_80_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ cpu.LCD0.row_2\[124\] cpu.LCD0.row_2\[116\] net1008 vssd1 vssd1 vccd1 vccd1
+ _01715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06765__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ net2109 net2214 net1007 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12398__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11604_ net2411 net241 net360 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ net1128 cpu.DM0.data_i\[6\] _06307_ _06345_ vssd1 vssd1 vccd1 vccd1 _06346_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14323_ clknet_leaf_57_clk _01436_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ cpu.RF0.registers\[16\]\[1\] net254 net369 vssd1 vssd1 vccd1 vccd1 _00953_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13814__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11610__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07596__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14254_ clknet_leaf_0_clk _01367_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ net2852 net128 net378 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14490__Q cpu.LCD0.row_2\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06931__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ clknet_leaf_19_clk _00385_ net1176 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10417_ _01812_ net269 _05626_ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08223__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14185_ clknet_leaf_105_clk _01298_ net1151 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11397_ net2636 net146 net388 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10030__B1 cpu.IM0.address_IM\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ clknet_leaf_48_clk _00316_ net1362 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[100\]
+ sky130_fd_sc_hd__dfstp_1
X_10348_ cpu.f0.i\[26\] _05577_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__nand2_1
XANTENNA__10581__A1 _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ clknet_leaf_53_clk _00247_ net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10279_ net1891 net728 _05523_ _05524_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__a22o_1
X_12018_ net1606 net165 net310 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__mux2_1
XANTENNA__07762__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11057__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13969_ clknet_leaf_76_clk _01082_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06510_ cpu.f0.num\[1\] cpu.f0.i\[1\] vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__or2_1
XANTENNA__10097__B1 cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07490_ cpu.RF0.registers\[1\]\[5\] net589 net584 cpu.RF0.registers\[2\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a22o_1
XANTENNA__06675__A a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13344__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06441_ cpu.CU0.opcode\[4\] cpu.CU0.opcode\[6\] _01847_ vssd1 vssd1 vccd1 vccd1 _01849_
+ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_17_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ cpu.CU0.funct3\[1\] _02108_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__nor2_1
X_06372_ a1.READ_I vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08111_ cpu.IM0.address_IM\[22\] net551 _03400_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_
+ sky130_fd_sc_hd__a22o_4
X_09091_ net305 _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__nor2_2
XANTENNA__07002__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11520__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ net668 _03323_ _03328_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__or4_2
XANTENNA_clkload43_A clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 _01690_ vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold912 cpu.RF0.registers\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 cpu.RF0.registers\[13\]\[6\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08214__B1 _03503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold934 cpu.LCD0.row_2\[91\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold945 cpu.LCD0.row_2\[48\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 cpu.RF0.registers\[6\]\[20\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 cpu.RF0.registers\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 cpu.RF0.registers\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10572__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09993_ _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__nor2_1
Xhold989 cpu.RF0.registers\[29\]\[26\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06776__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ cpu.RF0.registers\[9\]\[27\] net699 _04217_ _04219_ _04223_ vssd1 vssd1 vccd1
+ vccd1 _04235_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1013_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08768__C _02038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07672__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ net1080 cpu.RF0.registers\[25\]\[17\] net862 vssd1 vssd1 vccd1 vccd1 _04166_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout473_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ net522 _03115_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07740__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_A _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ net1042 cpu.RF0.registers\[31\]\[21\] net827 vssd1 vssd1 vccd1 vccd1 _03048_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout738_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06708_ cpu.CU0.opcode\[4\] cpu.CU0.opcode\[6\] cpu.CU0.opcode\[5\] vssd1 vssd1 vccd1
+ vccd1 _01999_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ cpu.RF0.registers\[2\]\[16\] net584 _02949_ _02955_ _02970_ vssd1 vssd1 vccd1
+ vccd1 _02979_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_36_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13248__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ _04163_ _04664_ _04201_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ a1.CPU_DAT_O\[7\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[7\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_97_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout905_A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1268_X net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13837__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ net452 _04569_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08309_ net442 _03597_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ _04278_ _04578_ _04286_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11430__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ net2443 net191 net394 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13987__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ net2587 net174 net404 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09548__A3 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__C1 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__A2 _01872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10202_ cpu.IM0.address_IM\[29\] _05443_ cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1
+ vccd1 _05465_ sky130_fd_sc_hd__a21o_1
X_11182_ net2548 net209 net411 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__mux2_1
XANTENNA__12812__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13217__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ net718 net135 _05401_ net631 vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__a31o_1
XANTENNA__12114__X _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _05324_ _05329_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nand2_1
XANTENNA__07582__C net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__B _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_0_clk _00936_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14612__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ clknet_leaf_93_clk _00867_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11815__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ net991 cpu.f0.write_data\[12\] vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ net2149 cpu.LCD0.row_2\[99\] net1002 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XANTENNA__14485__Q cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06926__C net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13685_ clknet_leaf_69_clk _00798_ net1328 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10897_ net1765 net170 net433 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ net2531 cpu.LCD0.row_2\[30\] net1005 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12567_ _01890_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__or2_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11340__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14306_ clknet_leaf_95_clk _01419_ net1215 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ net1864 net192 net370 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__mux2_1
X_12498_ _05521_ _06268_ _06281_ net262 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__o211a_1
XANTENNA__07757__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold208 cpu.DM0.readdata\[14\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 cpu.RF0.registers\[29\]\[3\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ clknet_leaf_88_clk _01350_ net1294 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11449_ net2425 net194 net379 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14168_ clknet_leaf_6_clk _01281_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ clknet_leaf_53_clk _00299_ net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[83\]
+ sky130_fd_sc_hd__dfrtp_1
X_14099_ clknet_leaf_67_clk _01212_ net1297 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ net1034 cpu.RF0.registers\[20\]\[23\] net780 vssd1 vssd1 vccd1 vccd1 _02281_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09046__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08588__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1270 net1272 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11863__X _05939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08660_ _03938_ _03942_ _03946_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or4_1
Xfanout1281 net1283 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1292 net1294 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08885__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ net543 _02869_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__or2_2
X_08591_ net948 cpu.RF0.registers\[8\]\[4\] net871 vssd1 vssd1 vccd1 vccd1 _03882_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11515__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07542_ cpu.IG0.Instr\[28\] net521 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09475__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07473_ net1060 cpu.RF0.registers\[23\]\[5\] net818 vssd1 vssd1 vccd1 vccd1 _02764_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08683__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07788__X _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ _04501_ _04502_ net453 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__mux2_1
X_06424_ cpu.c0.count\[9\] _01835_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12884__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06355_ cpu.LCD0.nextState\[3\] vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__inv_2
X_09143_ _04430_ _04433_ net456 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11250__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09074_ _04158_ net439 net466 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux2_1
XANTENNA__07643__D1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08125__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08025_ net947 cpu.RF0.registers\[10\]\[24\] net861 vssd1 vssd1 vccd1 vccd1 _03316_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1130_A a1.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 cpu.LCD0.row_2\[62\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold731 cpu.RF0.registers\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 cpu.RF0.registers\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 cpu.RF0.registers\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 cpu.RF0.registers\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 cpu.RF0.registers\[16\]\[28\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 cpu.RF0.registers\[30\]\[29\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 cpu.RF0.registers\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10390__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _05253_ _05257_ net629 _04792_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net938 cpu.RF0.registers\[15\]\[27\] net859 vssd1 vssd1 vccd1 vccd1 _04218_
+ sky130_fd_sc_hd__and3_1
XANTENNA__14635__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A _02035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1420 cpu.RF0.registers\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09163__A1 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1431 cpu.RF0.registers\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 net2837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 cpu.RF0.registers\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_24_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08858_ cpu.RF0.registers\[8\]\[16\] net708 net684 cpu.RF0.registers\[24\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__a22o_1
Xhold1453 cpu.RF0.registers\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 cpu.f0.data_adr\[9\] vssd1 vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 cpu.f0.data_adr\[22\] vssd1 vssd1 vccd1 vccd1 net2881 sky130_fd_sc_hd__dlygate4sd3_1
X_07809_ net1031 cpu.RF0.registers\[16\]\[22\] net831 vssd1 vssd1 vccd1 vccd1 _03100_
+ sky130_fd_sc_hd__and3_1
Xhold1486 cpu.RF0.registers\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net2892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 cpu.DM0.data_i\[24\] vssd1 vssd1 vccd1 vccd1 net2903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ cpu.RF0.registers\[8\]\[18\] net707 net695 cpu.RF0.registers\[17\]\[18\]
+ _04060_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1385_X net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ cpu.f0.data_adr\[31\] _04447_ net989 vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12818__Q cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ cpu.f0.data_adr\[11\] _04792_ net992 vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__mux2_1
XANTENNA__08674__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ clknet_leaf_86_clk _00583_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net2679 cpu.LCD0.row_1\[96\] net910 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XANTENNA__09218__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14015__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ cpu.DM0.readdata\[18\] net731 net500 _06234_ vssd1 vssd1 vccd1 vccd1 _01534_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08426__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06762__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11160__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12773__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14288__RESET_B net1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ net1408 _06217_ _06218_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10784__A1 cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ net2142 net239 net396 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ cpu.LCD0.row_2\[39\] _06004_ _06006_ cpu.LCD0.row_1\[39\] _06176_ vssd1 vssd1
+ vccd1 vccd1 _06177_ sky130_fd_sc_hd__a221o_1
XANTENNA__14165__CLK clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ clknet_leaf_6_clk _01135_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11234_ net1568 net131 net406 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10536__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__C1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ net2879 net146 net416 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__mux2_1
X_10116_ net715 net132 _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a21oi_1
X_11096_ net2848 net158 net422 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_42_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10047_ net626 _04734_ net1023 vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__o21a_1
Xhold80 _00173_ vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold91 _00168_ vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13806_ clknet_leaf_1_clk _00919_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09457__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ net2700 net252 net313 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__mux2_1
X_13737_ clknet_leaf_2_clk _00850_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10949_ cpu.CU0.funct3\[0\] _01848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10472__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13668_ clknet_leaf_96_clk _00781_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ cpu.LCD0.row_2\[21\] cpu.LCD0.row_2\[13\] net1000 vssd1 vssd1 vccd1 vccd1
+ _01612_ sky130_fd_sc_hd__mux2_1
XANTENNA__08417__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06672__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ clknet_leaf_105_clk _00712_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14508__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10224__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12764__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10775__A1 a1.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09917__B1 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10922__B _04601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _04734_ _05096_ _05119_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
XFILLER_0_10_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09761_ _03995_ _03996_ _04026_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__a21oi_1
X_14669__1391 vssd1 vssd1 vccd1 vccd1 _14669__1391/HI net1391 sky130_fd_sc_hd__conb_1
X_06973_ cpu.RF0.registers\[15\]\[25\] net590 net565 cpu.RF0.registers\[30\]\[25\]
+ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08712_ cpu.RF0.registers\[4\]\[0\] net678 net669 cpu.RF0.registers\[22\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a22o_1
X_09692_ _04964_ _04982_ _04981_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a21o_1
XANTENNA__09696__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _03931_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__and2_1
XANTENNA__07950__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout171_A _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06847__B net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08574_ cpu.RF0.registers\[0\]\[5\] net664 net550 vssd1 vssd1 vccd1 vccd1 _03865_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14038__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ cpu.RF0.registers\[3\]\[6\] net610 net608 cpu.RF0.registers\[24\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09853__C1 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07959__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ cpu.RF0.registers\[5\]\[1\] net602 _02732_ _02737_ _02738_ vssd1 vssd1 vccd1
+ vccd1 _02747_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06863__A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__X _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06407_ _01822_ _01823_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[1\] sky130_fd_sc_hd__and2_1
XFILLER_0_88_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13062__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07387_ _02669_ _02670_ _02671_ _02677_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout603_A _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14188__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12755__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ net462 net442 _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07397__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ cpu.RF0.registers\[3\]\[31\] net609 _04324_ _04327_ _04341_ vssd1 vssd1 vccd1
+ vccd1 _04348_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ cpu.RF0.registers\[0\]\[28\] net664 net550 vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__10518__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold550 cpu.RF0.registers\[19\]\[28\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 cpu.RF0.registers\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 cpu.f0.num\[18\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold583 cpu.RF0.registers\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1300_X net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 cpu.RF0.registers\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ cpu.IM0.address_IM\[10\] cpu.IM0.address_IM\[9\] _05219_ vssd1 vssd1 vccd1
+ vccd1 _05242_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ clknet_leaf_44_clk net1557 net1306 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07147__B1 cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 cpu.RF0.registers\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 cpu.RF0.registers\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ net2833 net178 net323 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
Xhold1272 cpu.RF0.registers\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1283 cpu.RF0.registers\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 cpu.RF0.registers\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11155__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14640_ clknet_leaf_31_clk _01741_ net1206 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09133__B _03698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ net1813 net168 net330 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XANTENNA__09439__A2 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10803_ net1692 net560 net539 _05749_ vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__a22o_1
X_14571_ clknet_leaf_61_clk net2484 net1345 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12443__A1 cpu.DM0.readdata\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ net2259 net185 net340 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_52_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13405__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08111__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10454__B1 _05640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13522_ clknet_leaf_60_clk _00635_ net1345 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ cpu.f0.data_adr\[6\] _04896_ net993 vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06773__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13453_ clknet_leaf_103_clk _00566_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10665_ net2600 cpu.LCD0.row_1\[79\] net903 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12404_ net1881 net733 _06225_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__o21a_1
XANTENNA__10206__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ clknet_leaf_84_clk _00497_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ cpu.LCD0.row_1\[2\] net2461 net898 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13555__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ cpu.LCD0.cnt_20ms\[11\] _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ cpu.LCD0.row_2\[94\] _05983_ _06007_ cpu.LCD0.row_2\[118\] _06160_ vssd1
+ vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ clknet_leaf_68_clk _01118_ net1324 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11217_ net2490 net194 net408 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_12197_ cpu.LCD0.row_2\[59\] _06000_ _06034_ cpu.LCD0.row_2\[27\] _06094_ vssd1 vssd1
+ vccd1 vccd1 _06095_ sky130_fd_sc_hd__a221o_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
X_11148_ net2090 net202 net416 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XANTENNA__09127__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ net1790 net218 net422 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XANTENNA__12131__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06667__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13085__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08102__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07310_ _02587_ _02588_ _02590_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__or4_2
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08290_ cpu.RF0.registers\[9\]\[13\] net701 net648 cpu.RF0.registers\[25\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a22o_1
XANTENNA__06683__A a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10996__A1 _03077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14139__RESET_B net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ net959 cpu.RF0.registers\[2\]\[9\] net769 vssd1 vssd1 vccd1 vccd1 _02532_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12198__B1 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__D net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07172_ cpu.RF0.registers\[7\]\[11\] net595 _02440_ _02443_ _02445_ vssd1 vssd1 vccd1
+ vccd1 _02463_ sky130_fd_sc_hd__a2111o_1
XANTENNA_wire773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09602__A2 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14480__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__A1 cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12922__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 _02605_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 _05942_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12370__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 _05939_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_6
X_09813_ _04497_ _04853_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__o21ai_1
Xfanout337 _05937_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_8
Xfanout359 _05931_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout386_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _04975_ _05034_ _04475_ _04903_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06956_ cpu.RF0.registers\[0\]\[26\] net617 _02243_ _02246_ vssd1 vssd1 vccd1 vccd1
+ _02247_ sky130_fd_sc_hd__o22a_2
XANTENNA__07129__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12579__B _06337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__B1 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _02794_ _03866_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__or2_1
X_06887_ net1038 cpu.RF0.registers\[16\]\[27\] net831 vssd1 vssd1 vccd1 vccd1 _02178_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1295_A net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13428__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08626_ cpu.RF0.registers\[17\]\[3\] net695 net658 cpu.RF0.registers\[13\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_A _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net950 cpu.RF0.registers\[4\]\[5\] net876 vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08629__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A1 cpu.DM0.readdata\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout818_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ net1057 cpu.RF0.registers\[29\]\[6\] net794 vssd1 vssd1 vccd1 vccd1 _02799_
+ sky130_fd_sc_hd__and3_1
X_08488_ net1106 cpu.RF0.registers\[26\]\[7\] net861 vssd1 vssd1 vccd1 vccd1 _03779_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13578__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07439_ net978 cpu.RF0.registers\[9\]\[1\] net760 vssd1 vssd1 vccd1 vccd1 _02730_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07852__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__B1 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12728__A2 cpu.DM0.dhit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ net30 net753 net563 net2813 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_21_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10739__B2 cpu.IM0.address_IM\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09109_ _02094_ _04379_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or2_1
XANTENNA__08016__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ net1127 _05608_ net267 net2547 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_21_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12120_ _05981_ net743 _05993_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__and3_4
XFILLER_0_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07080__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__Q cpu.IM0.address_IM\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ cpu.LCD0.cnt_500hz\[4\] _01955_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 cpu.RF0.registers\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 cpu.RF0.registers\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net273 _05886_ _05887_ net925 a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1
+ _00430_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_70_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14203__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
Xfanout871 net873 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
Xfanout882 net884 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_4
Xfanout893 net895 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_2
XANTENNA__06768__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__C net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ clknet_leaf_20_clk _00142_ net1169 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1080 cpu.RF0.registers\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 cpu.LCD0.row_2\[22\] vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net2602 net224 net324 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XANTENNA__14353__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12884_ clknet_leaf_1_clk cpu.c0.next_count\[15\] net1139 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ clknet_leaf_30_clk _01724_ net1207 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_83_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11835_ net1988 net243 net332 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12709__S net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11613__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ clknet_leaf_50_clk net2525 net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ net1801 net255 net341 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__mux2_1
XANTENNA__10737__B _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14493__Q cpu.LCD0.row_2\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06934__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ clknet_leaf_63_clk _00618_ net1343 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net991 _05005_ net287 net1016 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1
+ _05689_ sky130_fd_sc_hd__a32o_1
X_14485_ clknet_leaf_41_clk _01588_ net1257 vssd1 vssd1 vccd1 vccd1 cpu.IM0.address_IM\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11697_ net1701 net128 net350 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
X_14668__1390 vssd1 vssd1 vccd1 vccd1 _14668__1390/HI net1390 sky130_fd_sc_hd__conb_1
XANTENNA__12945__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13436_ clknet_leaf_12_clk _00549_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10648_ net2934 cpu.LCD0.row_1\[62\] net907 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__mux2_1
XANTENNA__06790__X _02081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08399__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13367_ clknet_leaf_65_clk _00480_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10579_ cpu.f0.write_data\[2\] _02679_ net995 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ cpu.LCD0.cnt_20ms\[3\] _05945_ net2926 vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a21o_1
X_13298_ clknet_leaf_34_clk cpu.RU0.next_FetchedData\[5\] net1248 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07765__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12249_ cpu.LCD0.row_2\[21\] _06003_ _06034_ cpu.LCD0.row_2\[29\] vssd1 vssd1 vccd1
+ vccd1 _06145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10899__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10902__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _01999_ _02082_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__nand2_2
XANTENNA__08571__A2 _02014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09325__Y _04616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ _03044_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2_1
XANTENNA__12104__B1 _06004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09054__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ net1081 cpu.RF0.registers\[24\]\[30\] net870 vssd1 vssd1 vccd1 vccd1 _02032_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08323__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net272 _04744_ _04750_ _04566_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_17_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06672_ a1.CPU_DAT_O\[8\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[8\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ net1078 cpu.RF0.registers\[31\]\[9\] net859 vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__and3_1
X_09391_ _04496_ _04672_ _04679_ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a211o_2
XANTENNA__07005__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09647__A_N net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11523__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ _03629_ _03631_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_47_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09284__B1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07429__A4 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload73_A clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08273_ cpu.IM0.address_IM\[15\] net554 _03562_ _03563_ vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13870__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ net956 cpu.RF0.registers\[15\]\[9\] net825 vssd1 vssd1 vccd1 vccd1 _02515_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07155_ net1043 cpu.RF0.registers\[24\]\[11\] net812 vssd1 vssd1 vccd1 vccd1 _02446_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_93_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12591__A0 cpu.IM0.address_IM\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__B net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13100__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ _02373_ _02374_ _02375_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__or4_1
XANTENNA__07675__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14226__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__B2 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1308_A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 _05839_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout156 net158 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout167 net168 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13250__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14376__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net180 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
X_07988_ net1092 cpu.RF0.registers\[30\]\[28\] net839 vssd1 vssd1 vccd1 vccd1 _03279_
+ sky130_fd_sc_hd__and3_1
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
XANTENNA__07770__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ _04029_ _04030_ _05017_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06939_ net954 cpu.RF0.registers\[9\]\[26\] net756 vssd1 vssd1 vccd1 vccd1 _02230_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _04946_ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_54_clk_X clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10121__A2 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ net492 _02760_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ net494 _04865_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ net2290 net181 net360 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
XANTENNA__10557__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12826__Q cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ net2286 net191 net366 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__mux2_1
XANTENNA__07825__A1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_X clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ net1500 net917 net751 a1.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 _00175_
+ sky130_fd_sc_hd__a22o_1
X_14270_ clknet_leaf_83_clk _01383_ net1273 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11482_ net2520 net196 net376 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
X_13221_ clknet_leaf_84_clk _00401_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10433_ net1125 _05634_ net264 net2097 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12117__X _06018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06770__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13152_ clknet_leaf_48_clk _00332_ net1361 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[116\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_76_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07053__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ cpu.f0.i\[28\] _05589_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07585__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12103_ _05981_ _05982_ _05995_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_72_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ clknet_leaf_53_clk _00263_ net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ cpu.f0.i\[17\] net541 _05526_ cpu.f0.i\[18\] vssd1 vssd1 vccd1 vccd1 _05538_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07882__A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ cpu.LCD0.cnt_20ms\[5\] _05948_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__and2_1
XANTENNA__10345__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _02028_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06929__C net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13985_ clknet_leaf_70_clk _01098_ net1298 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12936_ clknet_leaf_29_clk _00125_ net1202 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14413__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12867_ clknet_leaf_27_clk _00085_ net1183 vssd1 vssd1 vccd1 vccd1 a1.BUSY_O sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11343__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14606_ clknet_leaf_47_clk _01708_ net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[117\]
+ sky130_fd_sc_hd__dfstp_1
X_11818_ net1849 net183 net337 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
X_12798_ net2817 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__clkbuf_1
X_14537_ clknet_leaf_49_clk _01639_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09040__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net1980 net191 net342 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09281__A3 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14468_ clknet_leaf_22_clk _01578_ net1174 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14249__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ clknet_leaf_89_clk _00532_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_14399_ clknet_leaf_21_clk _01510_ net1178 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06680__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07044__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09991__B cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13273__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ net1077 cpu.RF0.registers\[25\]\[26\] net862 vssd1 vssd1 vccd1 vccd1 _04251_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__14399__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07911_ net957 cpu.RF0.registers\[8\]\[30\] net811 vssd1 vssd1 vccd1 vccd1 _03202_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07792__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08891_ cpu.RF0.registers\[31\]\[17\] net687 net677 cpu.RF0.registers\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11518__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07842_ cpu.RF0.registers\[4\]\[24\] net587 net574 cpu.RF0.registers\[9\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06555__A1 cpu.f0.state\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14398__Q cpu.IG0.Instr\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ net967 cpu.RF0.registers\[9\]\[21\] net757 vssd1 vssd1 vccd1 vccd1 _03064_
+ sky130_fd_sc_hd__and3_1
X_09512_ _02903_ _03630_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nor2_1
X_06724_ net936 cpu.RF0.registers\[8\]\[30\] net870 vssd1 vssd1 vccd1 vccd1 _02015_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09512__A _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net493 _04717_ _04718_ _04731_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a311o_4
X_06655_ net1712 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[23\] sky130_fd_sc_hd__and2_1
XANTENNA_fanout251_A _05774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06855__B net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11253__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09374_ _04163_ _04200_ _04664_ _04198_ _04091_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a311oi_4
X_06586_ _01956_ _01958_ _01959_ _01960_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__or4_2
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ cpu.RF0.registers\[9\]\[12\] net699 net638 cpu.RF0.registers\[26\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10811__A0 cpu.f0.data_adr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08256_ cpu.RF0.registers\[15\]\[15\] net683 _03541_ _03546_ vssd1 vssd1 vccd1 vccd1
+ _03547_ sky130_fd_sc_hd__a211o_1
XANTENNA__07283__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06871__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ cpu.RF0.registers\[13\]\[10\] net597 _02481_ _02487_ _02489_ vssd1 vssd1
+ vccd1 vccd1 _02498_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ net939 cpu.RF0.registers\[1\]\[21\] net883 vssd1 vssd1 vccd1 vccd1 _03478_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ cpu.RF0.registers\[14\]\[15\] net575 net565 cpu.RF0.registers\[30\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07069_ net974 cpu.RF0.registers\[11\]\[18\] net777 vssd1 vssd1 vccd1 vccd1 _02360_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _05346_ _05351_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11428__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_100_clk _00883_ net1213 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09496__B1 _04402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _03018_ net532 vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ net1578 cpu.LCD0.row_2\[115\] net1002 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__C net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11163__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net2299 net2233 net1005 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__mux2_1
XANTENNA__09141__B _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13146__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ net2287 net248 net360 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
XANTENNA__12398__A3 _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12583_ _01873_ _06334_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__nor2_2
XANTENNA__13877__RESET_B net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ clknet_leaf_57_clk _01435_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10802__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11534_ net1810 net236 net368 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ clknet_leaf_105_clk _01366_ net1156 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_49_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13296__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11465_ net1731 net136 net378 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14541__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ clknet_leaf_64_clk _00384_ net1307 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net1126 _01813_ net265 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ clknet_leaf_99_clk _01297_ net1232 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11396_ net1917 net149 net389 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XANTENNA__10030__A1 cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ clknet_leaf_53_clk net2661 net1351 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_10347_ cpu.f0.i\[26\] _05577_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13066_ clknet_leaf_52_clk _00246_ net1380 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ cpu.f0.i\[15\] _05518_ net725 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__o21a_1
XANTENNA__10318__C1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11338__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ net1773 net168 net311 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__mux2_1
XANTENNA__09723__B2 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10333__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06537__B2 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09035__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ clknet_leaf_73_clk _01081_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10097__B2 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ clknet_leaf_27_clk _00108_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ clknet_leaf_89_clk _01012_ net1280 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06675__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06440_ cpu.CU0.opcode\[4\] cpu.CU0.opcode\[6\] _01847_ vssd1 vssd1 vccd1 vccd1 _01848_
+ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_17_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14071__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ a1.WRITE_I vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13639__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11801__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ cpu.RF0.registers\[0\]\[22\] net661 net547 vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09090_ _04379_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06473__B1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08041_ cpu.RF0.registers\[2\]\[24\] net655 _03329_ _03330_ _03331_ vssd1 vssd1 vccd1
+ vccd1 _03332_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold902 cpu.RF0.registers\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold913 cpu.FetchedInstr\[30\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08214__A1 cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13789__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 cpu.FetchedInstr\[23\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 _01682_ vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold946 cpu.LCD0.row_2\[72\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09962__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold957 cpu.RF0.registers\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 cpu.LCD0.row_2\[90\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ cpu.IM0.address_IM\[12\] _05254_ cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1
+ vccd1 _05272_ sky130_fd_sc_hd__a21oi_1
Xhold979 cpu.RF0.registers\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07973__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09066__X _04357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ cpu.RF0.registers\[2\]\[27\] net654 _04218_ _04224_ _04225_ vssd1 vssd1 vccd1
+ vccd1 _04234_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07953__C net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A _04392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08874_ _04162_ _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1006_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ net1068 net633 net519 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07756_ net1042 cpu.RF0.registers\[28\]\[21\] net766 vssd1 vssd1 vccd1 vccd1 _03047_
+ sky130_fd_sc_hd__and3_1
X_06707_ cpu.f0.state\[5\] _01871_ net528 vssd1 vssd1 vccd1 vccd1 cpu.f0.next_write_i
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14414__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ cpu.RF0.registers\[7\]\[16\] net596 _02951_ _02963_ _02966_ vssd1 vssd1 vccd1
+ vccd1 _02978_ sky130_fd_sc_hd__a2111o_1
X_09426_ _04163_ _04201_ _04664_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06638_ a1.CPU_DAT_O\[6\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[6\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_97_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09357_ _02274_ _03372_ _04645_ _04646_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a22o_1
X_06569_ cpu.RU0.state\[6\] net2761 net1130 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_dhit
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11711__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__inv_2
XANTENNA__14564__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__X _03436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _04278_ _04286_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__and3_1
XANTENNA__09650__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__B2 cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ cpu.RF0.registers\[10\]\[14\] net692 net675 cpu.RF0.registers\[6\]\[14\]
+ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07008__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net1971 net196 net404 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08024__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10201_ cpu.IM0.address_IM\[30\] cpu.IM0.address_IM\[29\] _05443_ vssd1 vssd1 vccd1
+ vccd1 _05464_ sky130_fd_sc_hd__and3_1
X_11181_ net2501 net201 net411 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__mux2_1
XANTENNA__10851__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07964__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08959__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ cpu.IM0.address_IM\[24\] _05387_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08321__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11158__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _05335_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__and2b_1
XANTENNA__12852__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11512__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10997__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12130__X _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09469__A0 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ clknet_leaf_86_clk _00935_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14094__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13753_ clknet_leaf_42_clk _00866_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10965_ _02901_ net516 _05852_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06495__B _01883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08141__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ net2473 net2247 net1001 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
X_13684_ clknet_leaf_69_clk _00797_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07495__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10896_ net723 _05343_ _05815_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a22o_1
X_12635_ cpu.LCD0.row_2\[37\] cpu.LCD0.row_2\[29\] net997 vssd1 vssd1 vccd1 vccd1
+ _01628_ sky130_fd_sc_hd__mux2_1
XANTENNA__07878__Y _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11621__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ _01869_ _06312_ _06309_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07247__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12240__A2 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07400__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ net2882 net205 net370 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
XANTENNA__13931__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14305_ clknet_leaf_64_clk _01418_ net1309 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12497_ _05521_ _06268_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold209 cpu.DM0.readdata\[13\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ clknet_leaf_11_clk _01349_ net1228 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ net2438 net199 net381 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14167_ clknet_leaf_64_clk _01280_ net1302 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ net2415 net214 net388 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
X_13118_ clknet_leaf_54_clk net2317 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07773__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ clknet_leaf_70_clk _01211_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__C1 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ clknet_leaf_45_clk _00229_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12161__D1 _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
Xfanout1271 net1272 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13311__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__clkbuf_2
Xfanout1293 net1294 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__clkbuf_4
X_07610_ cpu.RF0.registers\[0\]\[12\] net620 _02894_ _02900_ vssd1 vssd1 vccd1 vccd1
+ _02901_ sky130_fd_sc_hd__o22a_2
XFILLER_0_55_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08590_ net1100 cpu.RF0.registers\[26\]\[4\] _02025_ vssd1 vssd1 vccd1 vccd1 _03881_
+ sky130_fd_sc_hd__and3_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07541_ net304 _02760_ _02795_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__and4_4
XFILLER_0_92_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13461__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09997__A cpu.IM0.address_IM\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14587__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ net1060 cpu.RF0.registers\[21\]\[5\] net798 vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09880__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11019__A0 cpu.f0.write_data\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ _03402_ net443 net460 vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__mux2_1
X_06423_ cpu.c0.count\[6\] cpu.c0.count\[7\] cpu.c0.count\[8\] _01826_ vssd1 vssd1
+ vccd1 vccd1 _01835_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11531__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nor2_1
XANTENNA__12231__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07948__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _03236_ _04294_ _04362_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o21a_2
XFILLER_0_44_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10793__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06854__A_N net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08024_ net1097 cpu.RF0.registers\[19\]\[24\] net836 vssd1 vssd1 vccd1 vccd1 _03315_
+ sky130_fd_sc_hd__and3_1
XANTENNA_wire856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold710 cpu.RF0.registers\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _01653_ vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold732 cpu.RF0.registers\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold743 cpu.LCD0.row_2\[107\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 cpu.RF0.registers\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 cpu.RF0.registers\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 cpu.RF0.registers\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 a1.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08779__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ net717 net134 _05256_ net629 vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a31o_1
Xhold798 cpu.RF0.registers\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ net1083 cpu.RF0.registers\[23\]\[27\] net844 vssd1 vssd1 vccd1 vccd1 _04217_
+ sky130_fd_sc_hd__and3_1
Xhold1410 a1.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07980__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1421 cpu.f0.num\[29\] vssd1 vssd1 vccd1 vccd1 net2827 sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ cpu.RF0.registers\[7\]\[16\] net651 net665 vssd1 vssd1 vccd1 vccd1 _04148_
+ sky130_fd_sc_hd__a21o_1
Xhold1432 cpu.RF0.registers\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout750_A _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1443 cpu.RF0.registers\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net2849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1454 cpu.RF0.registers\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net2860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1465 cpu.RF0.registers\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net2871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07808_ net959 cpu.RF0.registers\[1\]\[22\] net805 vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__and3_1
Xhold1476 cpu.RF0.registers\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net2882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08788_ _04075_ _04076_ _04077_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__or4_1
Xhold1487 cpu.FetchedInstr\[18\] vssd1 vssd1 vccd1 vccd1 net2893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 cpu.RF0.registers\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net2904 sky130_fd_sc_hd__dlygate4sd3_1
X_07739_ cpu.RF0.registers\[27\]\[20\] net592 net589 cpu.RF0.registers\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ net2331 net560 net538 _05711_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ _02758_ _04698_ _04699_ _04480_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a22o_1
XANTENNA__08019__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ cpu.LCD0.row_1\[87\] net2488 net902 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12758__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ cpu.DM0.data_i\[18\] net535 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and2_1
XANTENNA__12222__A2 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08316__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10565__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__Q cpu.IM0.address_IM\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ net1408 _06217_ net1368 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10784__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ net503 _05910_ _05920_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__and3_4
XFILLER_0_65_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ cpu.LCD0.row_2\[55\] _06011_ _06027_ cpu.LCD0.row_2\[47\] vssd1 vssd1 vccd1
+ vccd1 _06176_ sky130_fd_sc_hd__a22o_1
X_14021_ clknet_leaf_8_clk _01134_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09926__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ net2102 net136 net406 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__mux2_1
XANTENNA__14257__RESET_B net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ net2675 net148 net417 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
XANTENNA__13334__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ _05383_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12289__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ net1841 net162 net424 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
XANTENNA__08986__A _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ net126 _05321_ _05318_ net627 vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a211o_1
Xhold70 _01711_ vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 net78 vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11616__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 cpu.f0.write_data\[9\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14496__Q cpu.LCD0.row_2\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06937__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13805_ clknet_leaf_104_clk _00918_ net1156 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ cpu.RF0.registers\[30\]\[1\] net254 net313 vssd1 vssd1 vccd1 vccd1 _01401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10948_ _01849_ _02095_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or2_1
X_13736_ clknet_leaf_99_clk _00849_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10472__B2 a1.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ clknet_leaf_78_clk _00780_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10879_ net2294 net195 net431 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11351__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12618_ cpu.LCD0.row_2\[20\] cpu.LCD0.row_2\[12\] net1002 vssd1 vssd1 vccd1 vccd1
+ _01611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07768__C net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ clknet_leaf_84_clk _00711_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10224__A1 cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12549_ cpu.K0.keyvalid cpu.f0.state\[5\] vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10775__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_1 _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09917__A1 cpu.IG0.Instr\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ clknet_leaf_90_clk _01332_ net1278 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07928__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout519 _02210_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _04409_ _04724_ _04732_ net292 _04696_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__o221a_2
X_06972_ cpu.RF0.registers\[2\]\[25\] net585 net566 cpu.RF0.registers\[11\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
XANTENNA__13827__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08711_ cpu.RF0.registers\[21\]\[0\] net647 net639 cpu.RF0.registers\[26\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a22o_1
X_09691_ net304 _03899_ _04967_ _02795_ _03866_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__o32ai_1
XANTENNA__11526__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_2
X_08642_ net492 _03932_ _03900_ net482 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12851__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ _03853_ _03858_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__or3_2
XANTENNA__13977__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08105__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07524_ net979 cpu.RF0.registers\[12\]\[6\] net768 vssd1 vssd1 vccd1 vccd1 _02815_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07459__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07455_ cpu.RF0.registers\[12\]\[1\] net572 _02724_ _02734_ _02736_ vssd1 vssd1 vccd1
+ vccd1 _02746_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10463__B2 a1.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A _05938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06863__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A cpu.IG0.Instr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ cpu.c0.count\[1\] cpu.c0.count\[0\] vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__or2_1
XANTENNA__07311__Y _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07386_ cpu.RF0.registers\[18\]\[2\] net579 _02647_ _02656_ net622 vssd1 vssd1 vccd1
+ vccd1 _02677_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07678__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07040__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ net467 _03629_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
XANTENNA__10215__A1 cpu.IM0.address_IM\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1338_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ cpu.RF0.registers\[11\]\[31\] net567 _04329_ _04334_ _04345_ vssd1 vssd1
+ vccd1 vccd1 _04347_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07975__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14602__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _03287_ _03289_ _03294_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__and4bb_1
Xhold540 cpu.RF0.registers\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold551 cpu.RF0.registers\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__A2 a1.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold562 cpu.RF0.registers\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14350__RESET_B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 cpu.RF0.registers\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 cpu.RF0.registers\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 cpu.RF0.registers\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09958_ _02004_ _05146_ _05239_ _05240_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__o211a_1
X_08909_ net439 _04196_ _04197_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__nand3_2
X_09889_ cpu.IM0.address_IM\[4\] cpu.IM0.address_IM\[3\] cpu.IM0.address_IM\[2\] vssd1
+ vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and3_1
XANTENNA__11436__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1240 cpu.RF0.registers\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 cpu.RF0.registers\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 cpu.RF0.registers\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ net1986 net154 net322 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
Xhold1273 cpu.LCD0.row_1\[88\] vssd1 vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 cpu.RF0.registers\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06757__C net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1295 cpu.RF0.registers\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
X_11851_ net2736 net181 net332 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10802_ net285 _05747_ _05748_ net1014 cpu.IM0.address_IM\[25\] vssd1 vssd1 vccd1
+ vccd1 _05749_ sky130_fd_sc_hd__a32o_1
X_14570_ clknet_leaf_50_clk _01672_ net1375 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ net2132 net189 net338 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ net1622 net559 net537 _05699_ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a22o_1
X_13521_ clknet_leaf_77_clk _00634_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10454__B2 a1.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06773__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14132__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13452_ clknet_leaf_80_clk _00565_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10664_ cpu.LCD0.row_1\[70\] net2582 net907 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07870__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08046__A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ cpu.DM0.data_i\[10\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10206__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10863__X _05793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ clknet_leaf_82_clk _00496_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10595_ cpu.LCD0.row_1\[1\] net2130 net908 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
XANTENNA__10757__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12334_ _06207_ net1340 _06206_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14282__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ cpu.LCD0.row_1\[110\] _06009_ _06015_ cpu.LCD0.row_1\[6\] vssd1 vssd1 vccd1
+ vccd1 _06160_ sky130_fd_sc_hd__a22o_1
XANTENNA__10509__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ clknet_leaf_71_clk _01117_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ net2009 net198 net406 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
X_12196_ cpu.LCD0.row_2\[67\] _05988_ _06025_ cpu.LCD0.row_1\[59\] vssd1 vssd1 vccd1
+ vccd1 _06094_ sky130_fd_sc_hd__a22o_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
X_11147_ net1587 net213 net416 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XANTENNA__12874__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11078_ net1721 net220 net424 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XANTENNA__11346__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ cpu.IM0.address_IM\[16\] cpu.IM0.address_IM\[15\] _05284_ vssd1 vssd1 vccd1
+ vccd1 _05306_ sky130_fd_sc_hd__and3_1
XANTENNA__07125__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09043__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08882__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__B2 a1.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__C1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_65_clk _00832_ net1281 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ net956 cpu.RF0.registers\[7\]\[9\] net816 vssd1 vssd1 vccd1 vccd1 _02531_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07861__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ cpu.RF0.registers\[5\]\[11\] net603 _02450_ _02452_ _02453_ vssd1 vssd1 vccd1
+ vccd1 _02462_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_87_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07795__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__X _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10207__A2_N _05469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout316 _05942_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_8
XANTENNA__12370__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__C net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__B2 cpu.CU0.funct3\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout327 _05939_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
X_09812_ _05100_ _05101_ _05102_ _05099_ _04916_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o32a_1
Xfanout338 _05936_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10381__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout349 _05934_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_4
XANTENNA__14005__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ net477 _04402_ net291 _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a211o_1
X_06955_ _02237_ _02238_ _02244_ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__or4_1
XANTENNA__07961__C net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A _01767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _04870_ _04963_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__or2_1
X_06886_ net1050 net832 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__and2_1
XANTENNA__10133__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07035__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ cpu.RF0.registers\[7\]\[3\] net653 _03903_ _03907_ _03911_ vssd1 vssd1 vccd1
+ vccd1 _03916_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14155__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1288_A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08556_ net950 cpu.RF0.registers\[6\]\[5\] net852 vssd1 vssd1 vccd1 vccd1 _03847_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06874__A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ cpu.RF0.registers\[0\]\[6\] net619 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08487_ net1106 cpu.RF0.registers\[27\]\[7\] net881 vssd1 vssd1 vccd1 vccd1 _03778_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout713_A _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06593__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07438_ net1055 cpu.RF0.registers\[31\]\[1\] net828 vssd1 vssd1 vccd1 vccd1 _02729_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07369_ net976 cpu.RF0.registers\[12\]\[2\] net767 vssd1 vssd1 vccd1 vccd1 _02660_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07201__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09108_ _02094_ _04379_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_21_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10380_ cpu.f0.i\[2\] net268 vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__nand2_1
XANTENNA__07604__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ net1025 cpu.RF0.registers\[24\]\[31\] net811 vssd1 vssd1 vccd1 vccd1 _04330_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ cpu.LCD0.cnt_500hz\[4\] _01955_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__or2_1
XANTENNA__12897__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 cpu.RF0.registers\[27\]\[19\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold381 cpu.f0.write_data\[7\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold392 cpu.RF0.registers\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08565__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ net985 cpu.f0.write_data\[22\] vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_70_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout850 _02041_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08967__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout861 _02025_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_6
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_2
Xfanout883 net884 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
XANTENNA__06768__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12952_ clknet_leaf_20_clk _00141_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 cpu.RF0.registers\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 cpu.RF0.registers\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 _01613_ vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ cpu.RF0.registers\[27\]\[6\] net228 net323 vssd1 vssd1 vccd1 vccd1 _01310_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12883_ clknet_leaf_1_clk cpu.c0.next_count\[14\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[14\] sky130_fd_sc_hd__dfrtp_1
X_14622_ clknet_leaf_33_clk _01723_ net1246 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_83_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net1697 net248 net333 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__A cpu.CU0.funct3\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14648__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ clknet_leaf_50_clk _01655_ net1381 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_11765_ net1540 net236 net340 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10716_ _01944_ _01949_ cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__o21a_2
X_13504_ clknet_leaf_5_clk _00617_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_14484_ clknet_leaf_29_clk net929 net1209 vssd1 vssd1 vccd1 vccd1 cpu.RU0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ net1638 net138 net350 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XANTENNA__07843__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10647_ cpu.LCD0.row_1\[53\] cpu.LCD0.row_1\[61\] net900 vssd1 vssd1 vccd1 vccd1
+ _00277_ sky130_fd_sc_hd__mux2_1
X_13435_ clknet_leaf_14_clk _00548_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ clknet_leaf_59_clk _00479_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10578_ _05676_ cpu.LCD0.row_1\[1\] net896 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14201__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ net1369 _05947_ _06197_ _05957_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a31o_1
X_13297_ clknet_leaf_34_clk cpu.RU0.next_FetchedData\[4\] net1248 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12248_ cpu.LCD0.row_2\[13\] _05998_ _06037_ cpu.LCD0.row_1\[77\] _06143_ vssd1 vssd1
+ vccd1 vccd1 _06144_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09038__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12179_ cpu.LCD0.row_1\[98\] _06024_ _06027_ cpu.LCD0.row_2\[42\] vssd1 vssd1 vccd1
+ vccd1 _06078_ sky130_fd_sc_hd__a22o_1
XANTENNA__10902__A2 _05131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08877__C net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06678__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13052__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14178__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06740_ net1087 net873 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06671_ a1.CPU_DAT_O\[7\] net890 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[7\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11804__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ net1082 cpu.RF0.registers\[19\]\[9\] net835 vssd1 vssd1 vccd1 vccd1 _03701_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ _02604_ _04680_ _04480_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__o21a_1
XANTENNA__12407__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06694__A a1.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ _03630_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11091__A1 _05822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07295__B1 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ cpu.RF0.registers\[0\]\[15\] net664 net550 vssd1 vssd1 vccd1 vccd1 _03563_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07834__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08117__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07223_ net1035 cpu.RF0.registers\[17\]\[9\] net804 vssd1 vssd1 vccd1 vccd1 _02514_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11599__X _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07154_ net1043 cpu.RF0.registers\[22\]\[11\] net801 vssd1 vssd1 vccd1 vccd1 _02445_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07956__C net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12932__Q a1.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07085_ cpu.RF0.registers\[13\]\[18\] net597 _02351_ _02362_ _02363_ vssd1 vssd1
+ vccd1 vccd1 _02376_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1036_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_A _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08547__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout135 _05147_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 _05839_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_2
Xfanout168 _05822_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
X_07987_ net1092 cpu.RF0.registers\[26\]\[28\] net860 vssd1 vssd1 vccd1 vccd1 _03278_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ _04029_ _04030_ net513 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__a21oi_1
X_06938_ net958 cpu.RF0.registers\[2\]\[26\] net770 vssd1 vssd1 vccd1 vccd1 _02229_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10106__B1 cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13545__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _02410_ _03534_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__xor2_1
X_06869_ net1055 net782 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout830_A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ cpu.IM0.address_IM\[4\] net553 _03897_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_
+ sky130_fd_sc_hd__a22o_2
X_09588_ _04574_ _04807_ _04866_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08539_ _03826_ _03827_ _03828_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13695__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11550_ net2271 net205 net366 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XANTENNA__06891__X _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07825__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10501_ net1544 net917 net751 a1.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 _00174_
+ sky130_fd_sc_hd__a22o_1
Xwire514 _02111_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08027__C net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ net1738 net198 net374 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13220_ clknet_leaf_78_clk _00400_ net1315 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11302__X _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__A2 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ cpu.f0.i\[28\] net268 vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__nand2_1
XANTENNA__10573__B net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12842__Q cpu.f0.data_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__B1 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ clknet_leaf_53_clk net2527 net1357 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10363_ cpu.f0.i\[28\] _05589_ net308 vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10593__A0 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08250__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _05989_ _05995_ net557 vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_72_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13082_ clknet_leaf_55_clk _00262_ net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ net1435 net724 _05533_ _05537_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_72_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__inv_2
XANTENNA__12133__X _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14320__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 _02036_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12098__B1 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net693 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13984_ clknet_leaf_8_clk _01097_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__A3 _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ clknet_leaf_29_clk _00124_ net1202 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14470__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11624__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12866_ clknet_leaf_32_clk net732 net1249 vssd1 vssd1 vccd1 vccd1 cpu.DM0.enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14605_ clknet_leaf_49_clk _01707_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[116\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06945__C net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ net1993 net172 net335 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__mux2_1
X_12797_ cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14536_ clknet_leaf_49_clk _01638_ net1374 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12270__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ net2099 net207 net342 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__mux2_1
XANTENNA__07816__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10820__A1 _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ clknet_leaf_22_clk _01577_ net1174 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ net1973 net199 net350 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ clknet_leaf_99_clk _00531_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14398_ clknet_leaf_21_clk _01509_ net1178 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13418__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ clknet_leaf_8_clk _00462_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10584__B1 _05679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08219__A_N net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08529__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ net957 cpu.RF0.registers\[13\]\[30\] net791 vssd1 vssd1 vccd1 vccd1 _03201_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08890_ _04178_ _04179_ _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_36_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07841_ cpu.RF0.registers\[6\]\[24\] _02175_ net576 cpu.RF0.registers\[14\]\[24\]
+ _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a221o_1
XANTENNA__13568__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07772_ net967 cpu.RF0.registers\[3\]\[21\] net821 vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__and3_1
X_09511_ _02903_ _03630_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and2_1
X_06723_ net939 net870 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_49_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11534__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 _03990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ net302 _04732_ _04479_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06654_ net2073 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ _04055_ _04056_ _04165_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a21o_2
X_06585_ cpu.LCD0.cnt_500hz\[5\] cpu.LCD0.cnt_500hz\[7\] cpu.LCD0.cnt_500hz\[6\] cpu.LCD0.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__or4b_1
XANTENNA__09257__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12970__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _05778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08324_ cpu.RF0.registers\[5\]\[12\] net704 net636 cpu.RF0.registers\[16\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12261__B1 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08255_ cpu.RF0.registers\[1\]\[15\] net713 net678 cpu.RF0.registers\[4\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout411_A _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__B net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ cpu.RF0.registers\[16\]\[10\] net582 _02478_ _02480_ _02492_ vssd1 vssd1
+ vccd1 vccd1 _02497_ sky130_fd_sc_hd__a2111o_1
X_08186_ _03474_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12564__B2 _06329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ cpu.RF0.registers\[19\]\[15\] net615 net595 cpu.RF0.registers\[7\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XANTENNA__10575__A0 cpu.f0.write_data\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1320_A net1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14343__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07983__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ net1053 cpu.RF0.registers\[25\]\[18\] net759 vssd1 vssd1 vccd1 vccd1 _02359_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11709__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14493__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12935__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _04998_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__nand2b_1
X_10981_ net273 _05871_ _05872_ net925 net1562 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a32o_1
XANTENNA__09496__A1 _03664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ net1534 cpu.LCD0.row_2\[114\] net1001 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08319__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12837__Q cpu.f0.data_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12651_ cpu.LCD0.row_2\[53\] cpu.LCD0.row_2\[45\] net997 vssd1 vssd1 vccd1 vccd1
+ _01644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ net2648 net249 net361 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XANTENNA__12252__B1 _06036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ _06344_ net1538 _06320_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09799__A2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10802__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14321_ clknet_leaf_57_clk _01434_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11533_ net505 _05906_ _05907_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_78_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08471__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ clknet_leaf_80_clk _01365_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11464_ net2091 net140 net379 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07596__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10415_ net1126 _05625_ net265 net2134 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__a2bb2o_1
X_13203_ clknet_leaf_59_clk _00383_ net1347 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10871__X _05799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ net2324 net156 net386 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__mux2_1
X_14183_ clknet_leaf_82_clk _01296_ net1291 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08223__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__A _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13134_ clknet_leaf_54_clk net2312 net1345 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ net1508 net726 _05581_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09971__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13710__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ clknet_leaf_45_clk _00245_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[29\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09156__Y _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net308 _05521_ _05522_ net527 vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a22o_1
X_12016_ net2904 net183 net313 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13860__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06796__X _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ clknet_leaf_87_clk _01080_ net1286 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11354__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ clknet_leaf_22_clk _00107_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ clknet_leaf_102_clk _01011_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14216__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ clknet_leaf_24_clk _00068_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09051__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06370_ net1023 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14519_ clknet_leaf_55_clk _01621_ net1366 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13240__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14366__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06473__A1 a1.WRITE_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08040_ cpu.RF0.registers\[15\]\[24\] net683 net652 cpu.RF0.registers\[7\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12808__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold903 cpu.RF0.registers\[23\]\[29\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 cpu.RF0.registers\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold925 a1.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 cpu.RF0.registers\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_53_clk_X clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 cpu.RF0.registers\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold958 cpu.RF0.registers\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ cpu.IM0.address_IM\[13\] cpu.IM0.address_IM\[12\] _05254_ vssd1 vssd1 vccd1
+ vccd1 _05271_ sky130_fd_sc_hd__and3_1
Xhold969 _01681_ vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06776__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload29_A clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12958__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ cpu.RF0.registers\[10\]\[27\] net693 _04214_ _04215_ _04221_ vssd1 vssd1
+ vccd1 vccd1 _04233_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08873_ _04159_ _04160_ _04161_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout194_A _05804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_X clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ cpu.RF0.registers\[0\]\[22\] net617 _03110_ _03114_ vssd1 vssd1 vccd1 vccd1
+ _03115_ sky130_fd_sc_hd__o22a_2
XFILLER_0_93_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09478__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ cpu.RF0.registers\[0\]\[21\] net620 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__or2_1
XANTENNA__09478__B2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A _05931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06866__B net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A _02756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ cpu.RU0.state\[0\] _01945_ _01946_ _00005_ vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_read_i
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07686_ cpu.RF0.registers\[28\]\[16\] net578 _02953_ _02960_ net621 vssd1 vssd1 vccd1
+ vccd1 _02977_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06637_ a1.CPU_DAT_O\[5\] net894 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[5\]
+ sky130_fd_sc_hd__and2_1
X_09425_ _04686_ _04705_ _04714_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__or3_1
XANTENNA__10956__X _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout626_A _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06568_ net1130 cpu.RU0.state\[4\] vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and2b_2
X_09356_ _02275_ _03372_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06882__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08307_ net442 _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09287_ _04212_ _04282_ _04284_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__o21ai_2
X_06499_ cpu.K0.code\[0\] _01888_ cpu.K0.code\[1\] vssd1 vssd1 vccd1 vccd1 _01889_
+ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ cpu.RF0.registers\[1\]\[14\] net713 net660 cpu.RF0.registers\[30\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout995_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13733__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ net949 cpu.RF0.registers\[8\]\[20\] net872 vssd1 vssd1 vccd1 vccd1 _03460_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08205__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ _05461_ _05462_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and2_1
X_11180_ net1896 net213 net413 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10851__B _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11439__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _05398_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor2_1
XANTENNA__13883__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09364__A1_N net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__A cpu.IG0.Instr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ cpu.IM0.address_IM\[19\] _02315_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14239__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ clknet_leaf_68_clk _00934_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09469__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11174__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13752_ clknet_leaf_6_clk _00865_ net1146 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ net276 _05859_ _05860_ net928 net1767 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12703_ net2396 net2394 net1011 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
X_13683_ clknet_leaf_67_clk _00796_ net1298 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13263__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ cpu.DM0.readdata\[19\] net735 net719 vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o21a_1
XANTENNA__11902__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14389__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12225__B1 _06027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ cpu.LCD0.row_2\[36\] cpu.LCD0.row_2\[28\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12565_ _06330_ cpu.SR1.char_in\[2\] _06320_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ clknet_leaf_4_clk _01417_ net1144 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11516_ net2606 net175 net372 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12496_ _01808_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ clknet_leaf_92_clk _01348_ net1241 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11447_ net2476 net208 net381 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ net2410 net218 net386 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__mux2_1
X_14166_ clknet_leaf_57_clk _01279_ net1365 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08512__A _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10554__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11349__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ clknet_leaf_51_clk _00297_ net1379 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[81\]
+ sky130_fd_sc_hd__dfrtp_1
X_10329_ net1019 cpu.f0.i\[23\] _05556_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__or3_2
X_14097_ clknet_leaf_76_clk _01210_ net1335 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__B1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ clknet_leaf_48_clk _00228_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09046__C net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1250 net1254 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_4
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__clkbuf_2
Xfanout1272 net1300 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_2
Xfanout1283 net1300 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__clkbuf_2
Xfanout1294 net1299 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_2
XANTENNA__08885__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11084__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06686__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _02582_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07471_ cpu.RF0.registers\[0\]\[5\] net618 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__or2_1
XANTENNA__09997__B _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__A1 _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08683__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06422_ _01827_ _01828_ _01834_ vssd1 vssd1 vccd1 vccd1 cpu.c0.next_count\[7\] sky130_fd_sc_hd__and3_1
X_09210_ net444 net440 net461 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__mux2_1
XANTENNA__12216__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07798__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07891__B1 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12767__A1 cpu.f0.write_data\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13756__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net467 _03833_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nor2_1
XANTENNA__12767__B2 cpu.f0.i\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12209__A _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08435__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09072_ _03236_ _04294_ _04362_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__nor3_2
X_08023_ net1097 cpu.RF0.registers\[29\]\[24\] net849 vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08125__C net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold700 cpu.RF0.registers\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A _05810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold711 cpu.RF0.registers\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 cpu.f0.num\[8\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold733 cpu.RF0.registers\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _01698_ vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09518__A _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 cpu.RF0.registers\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12940__Q a1.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 cpu.RF0.registers\[8\]\[2\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11259__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold777 cpu.RF0.registers\[4\]\[17\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 cpu.LCD0.row_2\[16\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _05254_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__or2_1
Xhold799 cpu.RF0.registers\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13136__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__X _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net938 cpu.RF0.registers\[5\]\[27\] net866 vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__and3_1
Xhold1400 cpu.RF0.registers\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 cpu.RF0.registers\[0\]\[24\] vssd1 vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 cpu.LCD0.row_2\[66\] vssd1 vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ cpu.RF0.registers\[15\]\[16\] net682 net642 cpu.RF0.registers\[3\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__a22o_1
Xhold1433 cpu.RF0.registers\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1444 cpu.RF0.registers\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net2850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 cpu.LCD0.cnt_20ms\[3\] vssd1 vssd1 vccd1 vccd1 net2861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 a1.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net2872 sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ net1031 cpu.RF0.registers\[25\]\[22\] net756 vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__and3_1
Xhold1477 cpu.FetchedInstr\[16\] vssd1 vssd1 vccd1 vccd1 net2883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1488 cpu.RF0.registers\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net2894 sky130_fd_sc_hd__dlygate4sd3_1
X_08787_ cpu.RF0.registers\[7\]\[18\] net652 net649 cpu.RF0.registers\[14\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08108__D1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1499 cpu.RF0.registers\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net2905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14531__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ cpu.RF0.registers\[28\]\[20\] net577 net568 cpu.RF0.registers\[25\]\[20\]
+ _03027_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09320__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09871__A1 cpu.IM0.address_IM\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ net953 cpu.RF0.registers\[13\]\[16\] net790 vssd1 vssd1 vccd1 vccd1 _02960_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11722__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ _04482_ _04484_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__nand2_1
X_10680_ net2696 cpu.LCD0.row_1\[94\] net907 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12758__B2 cpu.f0.i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ net478 _04629_ _04595_ _04475_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08426__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ _06217_ net1368 _06216_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ net2246 net131 net398 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
X_12281_ cpu.LCD0.row_2\[7\] _06016_ _06036_ cpu.LCD0.row_1\[23\] _06174_ vssd1 vssd1
+ vccd1 vccd1 _06175_ sky130_fd_sc_hd__a221o_1
X_11232_ net2642 net140 net408 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__mux2_1
X_14020_ clknet_leaf_96_clk _01133_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10536__A3 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ cpu.RF0.registers\[4\]\[26\] net155 net414 vssd1 vssd1 vccd1 vccd1 _00594_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09147__B _03931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10114_ _05371_ _05373_ _05369_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a21o_1
X_11094_ net2649 net179 net423 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
XANTENNA__14061__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12789__A cpu.RF0.registers\[0\]\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _05319_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__nor2_1
Xhold60 cpu.f0.write_data\[8\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 cpu.f0.write_data\[20\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 _00166_ vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net83 vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ clknet_leaf_87_clk _00917_ net1289 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11996_ net1717 net237 net312 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__mux2_1
XANTENNA__13779__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13735_ clknet_leaf_82_clk _00848_ net1288 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10947_ _01849_ _02095_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09610__B _04025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_11_clk _00779_ net1225 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08507__A _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ _05286_ _05803_ _02002_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__mux2_4
XFILLER_0_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12749__B2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12617_ cpu.LCD0.row_2\[19\] net2831 net997 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XANTENNA__13009__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ clknet_leaf_89_clk _00710_ net1280 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ _01870_ _06314_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__or3b_4
XFILLER_0_42_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12479_ net1021 cpu.f0.i\[8\] _06264_ cpu.f0.i\[9\] vssd1 vssd1 vccd1 vccd1 _06270_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_2 _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13159__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ clknet_leaf_100_clk _01331_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14404__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11079__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14149_ clknet_leaf_11_clk _01262_ net1222 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06971_ cpu.RF0.registers\[27\]\[25\] net591 _02260_ _02261_ vssd1 vssd1 vccd1 vccd1
+ _02262_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08710_ _03997_ _03998_ _03999_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__or4_1
XANTENNA__11807__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09690_ _04980_ _04870_ _03798_ _02582_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14554__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1080 net1082 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_2
X_08641_ net471 net468 net457 net482 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a31o_1
XANTENNA_wire809_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1091 net1109 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10160__A1 cpu.IM0.address_IM\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__A cpu.IM0.address_IM\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ _03859_ _03860_ _03861_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload96_A clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ net978 cpu.RF0.registers\[1\]\[6\] net807 vssd1 vssd1 vccd1 vccd1 _02814_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11542__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07454_ cpu.RF0.registers\[24\]\[1\] net608 _02723_ _02729_ _02742_ vssd1 vssd1 vccd1
+ vccd1 _02745_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07864__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07959__C net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06405_ cpu.c0.count\[1\] cpu.c0.count\[0\] vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07321__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07385_ _02672_ _02673_ _02674_ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__or4_2
XANTENNA__09605__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09055_ net1026 cpu.RF0.registers\[25\]\[31\] net756 vssd1 vssd1 vccd1 vccd1 _04346_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07092__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1233_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08006_ cpu.RF0.registers\[12\]\[28\] net697 net667 _03295_ _03296_ vssd1 vssd1 vccd1
+ vccd1 _03297_ sky130_fd_sc_hd__a2111oi_1
Xhold530 cpu.RF0.registers\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07694__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14084__CLK clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 cpu.RF0.registers\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 cpu.RF0.registers\[5\]\[22\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__A3 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 cpu.RF0.registers\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 cpu.RF0.registers\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 cpu.DM0.readdata\[27\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 a1.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _05235_ _05238_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08908_ net439 _04196_ _04197_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__and3_1
XANTENNA__14390__RESET_B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _02004_ _05146_ _05175_ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o211a_1
Xhold1230 cpu.RF0.registers\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1241 cpu.RF0.registers\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1252 cpu.RF0.registers\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ net1075 cpu.RF0.registers\[16\]\[16\] net841 vssd1 vssd1 vccd1 vccd1 _04130_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06400__A cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13921__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1263 cpu.RF0.registers\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _00312_ vssd1 vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1285 cpu.LCD0.row_2\[49\] vssd1 vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 cpu.RF0.registers\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ net1878 net170 net331 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ net986 cpu.f0.data_adr\[25\] vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or2_2
XANTENNA__08647__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net2025 net207 net338 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__mux2_1
XANTENNA__09844__B2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11452__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ clknet_leaf_75_clk _00633_ net1333 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07502__Y _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ net285 _05697_ _05698_ net1015 cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1
+ vccd1 _05699_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07231__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11024__Y _05902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13451_ clknet_leaf_90_clk _00564_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10663_ cpu.LCD0.row_1\[69\] cpu.LCD0.row_1\[77\] net900 vssd1 vssd1 vccd1 vccd1
+ _00293_ sky130_fd_sc_hd__mux2_1
X_12402_ net1436 net732 _06224_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__o21a_1
XANTENNA__12600__A0 cpu.LCD0.row_2\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ cpu.LCD0.row_1\[0\] net2457 net909 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13382_ clknet_leaf_7_clk _00495_ net1149 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13301__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14427__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12333_ cpu.LCD0.cnt_20ms\[10\] cpu.LCD0.cnt_20ms\[9\] _06203_ vssd1 vssd1 vccd1
+ vccd1 _06207_ sky130_fd_sc_hd__and3_1
XANTENNA__12136__X _06037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_12264_ cpu.LCD0.row_2\[22\] _06003_ _06022_ cpu.LCD0.row_2\[126\] _06158_ vssd1
+ vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ clknet_leaf_69_clk _01116_ net1325 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11215_ net1627 net209 net406 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
X_12195_ cpu.LCD0.row_2\[123\] _06022_ _06036_ cpu.LCD0.row_1\[19\] _06092_ vssd1
+ vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13451__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XANTENNA__14577__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__07386__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_11146_ net2885 net216 net414 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11627__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11077_ cpu.RF0.registers\[2\]\[7\] net226 net423 vssd1 vssd1 vccd1 vccd1 _00511_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07138__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__A2 _06030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10028_ _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__and2_1
XANTENNA__10142__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09621__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11979_ net1663 net206 net314 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11362__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_70_clk _00831_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ clknet_leaf_78_clk _00762_ net1319 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12198__A2 _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07170_ cpu.RF0.registers\[13\]\[11\] net597 _02448_ _02454_ _02455_ vssd1 vssd1
+ vccd1 vccd1 _02461_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_13_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09063__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06821__A1 cpu.CU0.funct3\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12206__B _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 _02604_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
Xfanout317 _05942_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_4
X_09811_ _04385_ _04688_ net278 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__o21ai_1
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_6
Xfanout339 _05936_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13944__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _04396_ net299 _04976_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__mux2_1
X_06954_ cpu.RF0.registers\[5\]\[26\] net603 _02217_ _02219_ _02234_ vssd1 vssd1 vccd1
+ vccd1 _02245_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07129__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__A2 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _04870_ _04963_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__nor2_1
XANTENNA__10133__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06885_ net962 cpu.RF0.registers\[6\]\[27\] net801 vssd1 vssd1 vccd1 vccd1 _02176_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout274_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ cpu.RF0.registers\[24\]\[3\] net685 net639 cpu.RF0.registers\[26\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a22o_1
XANTENNA__06862__B_N net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08555_ net1105 cpu.RF0.registers\[30\]\[5\] net840 vssd1 vssd1 vccd1 vccd1 _03846_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09826__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__B net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ cpu.IG0.Instr\[26\] net520 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__and2_2
XANTENNA__09250__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07837__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ net950 cpu.RF0.registers\[14\]\[7\] net839 vssd1 vssd1 vccd1 vccd1 _03777_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07301__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ net1056 cpu.RF0.registers\[18\]\[1\] net772 vssd1 vssd1 vccd1 vccd1 _02728_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1350_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__A2 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ net1054 cpu.RF0.registers\[16\]\[2\] net832 vssd1 vssd1 vccd1 vccd1 _02659_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10739__A3 _05703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ net438 _04358_ net295 vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_21_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08262__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07299_ cpu.RF0.registers\[3\]\[4\] net610 net581 cpu.RF0.registers\[16\]\[4\] _02589_
+ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a221o_1
X_09038_ net1028 cpu.RF0.registers\[19\]\[31\] net820 vssd1 vssd1 vccd1 vccd1 _04329_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__C net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 cpu.RF0.registers\[0\]\[22\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 cpu.RF0.registers\[5\]\[5\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 cpu.RF0.registers\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 cpu.RF0.registers\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net282 _05885_ net986 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09762__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _02052_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout851 net852 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_8
Xfanout862 net864 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09425__B _04705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 _02013_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09514__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout884 _02006_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout895 cpu.RU0.next_ihit vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_2
X_12951_ clknet_leaf_20_clk _00140_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 _01622_ vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1071 cpu.LCD0.row_1\[18\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net1659 net235 net324 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
Xhold1082 cpu.LCD0.row_1\[95\] vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 cpu.LCD0.row_2\[41\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ clknet_leaf_1_clk cpu.c0.next_count\[13\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[13\] sky130_fd_sc_hd__dfrtp_1
X_14621_ clknet_leaf_30_clk _01722_ net1245 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_83_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11833_ net2250 net250 net333 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11182__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11035__X _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A0 _03115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14552_ clknet_leaf_51_clk _01654_ net1373 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11764_ net506 _05765_ _05915_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__and3_4
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13503_ clknet_leaf_0_clk _00616_ net1138 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ net1013 cpu.RU0.state\[0\] net558 vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14483_ clknet_leaf_30_clk _00006_ net1208 vssd1 vssd1 vccd1 vccd1 cpu.RU0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ net2533 net142 net352 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XANTENNA__11910__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13817__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ clknet_leaf_96_clk _00547_ net1234 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ cpu.LCD0.row_1\[52\] cpu.LCD0.row_1\[60\] net904 vssd1 vssd1 vccd1 vccd1
+ _00276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ clknet_leaf_73_clk _00478_ net1337 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10577_ cpu.f0.write_data\[1\] _02754_ net995 vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12316_ cpu.LCD0.cnt_20ms\[3\] _05945_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__or2_1
XANTENNA__07461__D1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13296_ clknet_leaf_33_clk cpu.RU0.next_FetchedData\[3\] net1247 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[3\] sky130_fd_sc_hd__dfrtp_1
X_12247_ cpu.LCD0.row_2\[85\] _05990_ _06028_ cpu.LCD0.row_1\[117\] vssd1 vssd1 vccd1
+ vccd1 _06143_ sky130_fd_sc_hd__a22o_1
XANTENNA__09202__C1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14241__RESET_B net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A1 cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ cpu.LCD0.row_2\[82\] _05990_ _06030_ cpu.LCD0.row_1\[42\] _06076_ vssd1 vssd1
+ vccd1 vccd1 _06077_ sky130_fd_sc_hd__a221o_1
XANTENNA__08520__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11357__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11129_ net1791 net157 net418 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12042__A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__A0 _03594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__A2 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09054__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06670_ a1.CPU_DAT_O\[6\] net891 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedData\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_56_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13347__CLK clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07531__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__A1 _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06694__B net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08340_ _02903_ _03595_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07142__Y _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08271_ _03555_ _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__X _05736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13497__CLK clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11820__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07222_ net1036 cpu.RF0.registers\[29\]\[9\] net790 vssd1 vssd1 vccd1 vccd1 _02513_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ net966 cpu.RF0.registers\[14\]\[11\] net762 vssd1 vssd1 vccd1 vccd1 _02444_
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkload59_A clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__Y _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08795__A1 cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09992__B1 cpu.IM0.address_IM\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ cpu.RF0.registers\[15\]\[18\] net590 _02360_ _02361_ _02368_ vssd1 vssd1
+ vccd1 vccd1 _02375_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_93_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10960__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__B1 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06558__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 _05149_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_4
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 net139 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _05839_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout158 _05834_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14122__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 _05822_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
X_07986_ net1093 cpu.RF0.registers\[23\]\[28\] net845 vssd1 vssd1 vccd1 vccd1 _03277_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_96_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07770__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ net494 _05006_ _05012_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a211o_2
X_06937_ net954 cpu.RF0.registers\[10\]\[26\] net786 vssd1 vssd1 vccd1 vccd1 _02228_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10106__A1 cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _02410_ _03535_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__nor2_1
X_06868_ net1072 net1069 net1065 net1067 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__nor4b_1
XANTENNA__14272__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ cpu.RF0.registers\[0\]\[4\] net663 net549 vssd1 vssd1 vccd1 vccd1 _03898_
+ sky130_fd_sc_hd__o21a_1
X_09587_ _04441_ net272 net277 _04877_ _04871_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout823_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ cpu.CU0.opcode\[2\] cpu.CU0.opcode\[5\] cpu.CU0.opcode\[1\] cpu.CU0.opcode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ cpu.RF0.registers\[5\]\[6\] net704 _03805_ _03814_ _03816_ vssd1 vssd1 vccd1
+ vccd1 _03829_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ net1093 cpu.RF0.registers\[18\]\[8\] net854 vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11730__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ net1485 net922 net747 a1.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 _00173_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09027__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ net1981 net211 net374 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XANTENNA__12864__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ net1125 _05633_ net264 net2232 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08235__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__A3 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11031__A cpu.IG0.Instr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09983__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13150_ clknet_leaf_54_clk net2236 net1346 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10362_ net527 _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__nand2_1
XANTENNA__10593__A1 cpu.LCD0.row_1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ cpu.LCD0.row_2\[56\] _06000_ _06001_ cpu.LCD0.row_1\[64\] _05999_ vssd1 vssd1
+ vccd1 vccd1 _06002_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_72_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13081_ clknet_leaf_45_clk _00261_ net1353 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[45\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12561__S _06320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ net307 _05536_ net728 vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_72_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12032_ cpu.LCD0.cnt_20ms\[4\] cpu.LCD0.cnt_20ms\[3\] _05945_ vssd1 vssd1 vccd1 vccd1
+ _05948_ sky130_fd_sc_hd__and3_1
Xhold190 cpu.RF0.registers\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08340__A _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _02047_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_89_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout681 _02036_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout692 net693 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
X_13983_ clknet_leaf_0_clk _01096_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12797__A cpu.RF0.registers\[0\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11905__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ clknet_leaf_28_clk _00123_ net1189 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12865_ clknet_leaf_24_clk _00084_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14604_ clknet_leaf_46_clk _01706_ net1358 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_11816_ net2470 net185 net336 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12796_ net1766 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ clknet_leaf_55_clk net2234 net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_11747_ net2026 net173 net343 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__mux2_1
XANTENNA__08474__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11640__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ clknet_leaf_22_clk _01576_ net1174 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09018__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11678_ net1867 net208 net350 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ clknet_leaf_2_clk _00530_ net1157 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ cpu.LCD0.row_1\[35\] net2389 net899 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ clknet_leaf_21_clk _01508_ net1177 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ clknet_leaf_96_clk _00461_ net1230 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10584__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06788__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10780__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14145__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13279_ clknet_leaf_21_clk cpu.RU0.next_FetchedInstr\[18\] net1176 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09726__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10336__A1 cpu.f0.i\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11087__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06689__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ cpu.RF0.registers\[8\]\[24\] net612 net589 cpu.RF0.registers\[1\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14295__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ net1042 cpu.RF0.registers\[21\]\[21\] net796 vssd1 vssd1 vccd1 vccd1 _03062_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09510_ net277 _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nand2_1
XANTENNA__11815__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06722_ net1114 net1116 net1112 net1110 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_95_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08701__A1 cpu.IM0.address_IM\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ net479 _04651_ _04723_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_49_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06653_ net1825 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[21\] sky130_fd_sc_hd__and2_1
XFILLER_0_8_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ net511 _04642_ _04643_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o31a_2
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06584_ cpu.LCD0.cnt_500hz\[8\] cpu.LCD0.cnt_500hz\[13\] cpu.LCD0.cnt_500hz\[12\]
+ cpu.LCD0.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__or4b_1
XANTENNA__12887__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06562__A_N net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08128__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ cpu.RF0.registers\[1\]\[12\] net714 net642 cpu.RF0.registers\[3\]\[12\] _03613_
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07032__C net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout237_A _05770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11550__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08254_ cpu.RF0.registers\[20\]\[15\] net709 net639 cpu.RF0.registers\[26\]\[15\]
+ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12943__Q a1.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07205_ cpu.RF0.registers\[19\]\[10\] net615 net578 cpu.RF0.registers\[28\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a22o_1
XANTENNA__12013__A1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ _03472_ _03473_ net444 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout404_A _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07136_ cpu.RF0.registers\[24\]\[15\] net607 net597 cpu.RF0.registers\[13\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10575__A1 _02716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ net974 cpu.RF0.registers\[6\]\[18\] net802 vssd1 vssd1 vccd1 vccd1 _02358_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1313_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09256__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14638__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__A1 _05479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13512__CLK clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__B2 cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ cpu.RF0.registers\[4\]\[29\] net679 _03240_ _03247_ _03252_ vssd1 vssd1 vccd1
+ vccd1 _03260_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout940_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ net451 _03992_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__nand2_1
X_10980_ net985 cpu.f0.write_data\[16\] vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09496__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _02384_ net441 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ cpu.LCD0.row_2\[52\] cpu.LCD0.row_2\[44\] net1003 vssd1 vssd1 vccd1 vccd1
+ _01643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14018__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11601_ net1763 net255 net361 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _06308_ _06342_ _06343_ net1129 vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09799__A3 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11460__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ clknet_leaf_58_clk _01433_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ net2911 net129 net370 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ clknet_leaf_90_clk _01364_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11463_ net2364 net146 net379 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ clknet_leaf_74_clk _00382_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10414_ net1020 net269 vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__nand2_1
X_14182_ clknet_leaf_6_clk _01295_ net1147 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10566__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11394_ net2055 net162 net388 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13133_ clknet_leaf_52_clk net2509 net1378 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_10345_ net526 _05576_ _05577_ _05580_ net724 vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o311a_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09166__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ clknet_leaf_48_clk _00244_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_10276_ cpu.f0.i\[15\] _05521_ net540 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12015_ net1964 net170 net311 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10105__A cpu.IM0.address_IM\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07734__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11635__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13966_ clknet_leaf_2_clk _01079_ net1153 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12917_ clknet_leaf_25_clk _00106_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08695__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ clknet_leaf_104_clk _01010_ net1152 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09892__C1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ clknet_leaf_31_clk _00067_ net1200 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08447__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ net1551 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11370__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14518_ clknet_leaf_45_clk _01620_ net1310 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[29\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14449_ clknet_leaf_26_clk _01559_ net1185 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_90_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 cpu.RF0.registers\[7\]\[17\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13535__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold915 cpu.RF0.registers\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 cpu.RF0.registers\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold937 cpu.RF0.registers\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold948 cpu.RF0.registers\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold959 cpu.LCD0.row_1\[41\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ net715 net132 _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07973__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08941_ cpu.RF0.registers\[8\]\[27\] net708 _04213_ _04220_ _04222_ vssd1 vssd1 vccd1
+ vccd1 _04232_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12214__B _06111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08411__C net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _04160_ _04161_ _04159_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a21o_1
XANTENNA__13685__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__X _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _03105_ _03111_ _03112_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__or4_1
XANTENNA__07027__C net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__inv_2
XANTENNA__12938__Q a1.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ cpu.RU0.state\[0\] _01949_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__and2_1
X_07685_ _02972_ _02973_ _02974_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or4_1
XANTENNA__08686__B1 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout354_A _05932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1096_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09424_ _04686_ _04705_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__nor3_1
X_06636_ a1.CPU_DAT_O\[4\] net895 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[4\]
+ sky130_fd_sc_hd__and2_1
X_09355_ _02274_ net434 _04644_ net293 net288 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__o221a_1
X_06567_ net1130 cpu.RU0.state\[2\] vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_ihit sky130_fd_sc_hd__and2b_1
XFILLER_0_30_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06882__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ _02940_ _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09286_ net493 _04556_ _04557_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a31o_2
XFILLER_0_30_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10796__A1 a1.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06498_ cpu.K0.code\[3\] cpu.K0.code\[2\] vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07697__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_7_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__A2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10796__B2 _05744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ cpu.RF0.registers\[9\]\[14\] net700 net669 cpu.RF0.registers\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1469_A a1.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__X _05866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ cpu.RF0.registers\[7\]\[20\] net652 _03457_ _03458_ net668 vssd1 vssd1 vccd1
+ vccd1 _03459_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14460__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout988_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ net523 _02408_ _02409_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_43_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12902__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ cpu.RF0.registers\[15\]\[22\] net682 net654 cpu.RF0.registers\[2\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a22o_1
XANTENNA__07058__X _02349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ _05392_ _05395_ _05397_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08321__C net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10061_ cpu.IM0.address_IM\[19\] _02315_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__and2_1
XANTENNA__07218__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__B1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__A1 _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A _04911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__C1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__A1 a1.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11455__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ clknet_leaf_15_clk _00933_ net1242 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12848__Q cpu.f0.data_adr\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ clknet_leaf_64_clk _00864_ net1301 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10963_ net987 cpu.f0.write_data\[11\] vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_82_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13408__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ net2404 cpu.LCD0.row_2\[96\] net1010 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XANTENNA__08141__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10484__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13682_ clknet_leaf_60_clk _00795_ net1344 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ net737 _04683_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12633_ cpu.LCD0.row_2\[35\] net2559 net999 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11190__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12564_ net1128 cpu.DM0.data_i\[2\] _06307_ _06329_ vssd1 vssd1 vccd1 vccd1 _06330_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13558__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14303_ clknet_leaf_0_clk _01416_ net1143 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14014__RESET_B net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11515_ net2301 net195 net371 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__mux2_1
XANTENNA__07400__C net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__X _05807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ net262 _06279_ _06280_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ clknet_leaf_94_clk _01347_ net1236 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11446_ net2445 net201 net378 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14165_ clknet_leaf_74_clk _01278_ net1327 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11377_ net1920 net222 net388 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13116_ clknet_leaf_50_clk _00296_ net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10328_ net1018 _05560_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__xnor2_1
X_14096_ clknet_leaf_74_clk _01209_ net1320 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13047_ clknet_leaf_47_clk _00227_ net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ net526 _05506_ _05507_ net724 vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__o31a_1
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_2
Xfanout1251 net1254 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1262 net1267 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_2
Xfanout1273 net1275 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11365__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1284 net1287 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__clkbuf_4
Xfanout1295 net1299 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07144__A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08668__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ clknet_leaf_89_clk _01062_ net1292 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_73_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08132__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ cpu.IG0.Instr\[25\] net521 net544 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09880__A2 _05030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06421_ _01829_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__or2_1
XANTENNA__12216__A1 cpu.LCD0.row_1\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12767__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09140_ net462 _03797_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__nor2_1
XANTENNA__12209__B _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09071_ _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12925__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08022_ net947 cpu.RF0.registers\[1\]\[24\] net884 vssd1 vssd1 vccd1 vccd1 _03313_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_13_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload41_A clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 cpu.RF0.registers\[8\]\[10\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 cpu.RF0.registers\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 cpu.f0.num\[13\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08199__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold734 cpu.f0.num\[3\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 cpu.RF0.registers\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold756 cpu.RF0.registers\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 cpu.LCD0.row_2\[25\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 cpu.RF0.registers\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07319__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09973_ cpu.IM0.address_IM\[11\] _05242_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold789 _01607_ vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ net1084 cpu.RF0.registers\[29\]\[27\] net848 vssd1 vssd1 vccd1 vccd1 _04215_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13390__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1401 cpu.RF0.registers\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1412 cpu.K0.code\[3\] vssd1 vssd1 vccd1 vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ cpu.RF0.registers\[6\]\[16\] net674 net640 cpu.RF0.registers\[19\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a22o_1
Xhold1423 cpu.RF0.registers\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 cpu.RF0.registers\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1445 cpu.c0.count\[16\] vssd1 vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ net1032 cpu.RF0.registers\[30\]\[22\] net762 vssd1 vssd1 vccd1 vccd1 _03097_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1456 cpu.RF0.registers\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net2862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1467 cpu.RF0.registers\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net2873 sky130_fd_sc_hd__dlygate4sd3_1
X_08786_ cpu.RF0.registers\[27\]\[18\] net712 _02059_ cpu.RF0.registers\[25\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a22o_1
Xhold1478 cpu.RF0.registers\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net2884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 cpu.RF0.registers\[0\]\[20\] vssd1 vssd1 vccd1 vccd1 net2895 sky130_fd_sc_hd__dlygate4sd3_1
X_07737_ cpu.RF0.registers\[23\]\[20\] net613 net607 cpu.RF0.registers\[24\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ net953 cpu.RF0.registers\[4\]\[16\] net780 vssd1 vssd1 vccd1 vccd1 _02959_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_95_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__A2 _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ _02089_ _03300_ net437 _03268_ net453 net460 vssd1 vssd1 vccd1 vccd1 _04698_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__13700__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06619_ _01972_ _01974_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout903_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ cpu.RF0.registers\[4\]\[12\] net586 _02872_ _02881_ _02885_ vssd1 vssd1 vccd1
+ vccd1 _02890_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1266_X net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__A2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ _04462_ _04470_ net473 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08316__C net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ net445 net295 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__nand2_1
XANTENNA__07220__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ net1573 net138 net398 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
XANTENNA__13850__CLK clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12280_ cpu.LCD0.row_1\[55\] _06019_ _06024_ cpu.LCD0.row_1\[103\] vssd1 vssd1 vccd1
+ vccd1 _06174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08613__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11231_ net2837 net145 net407 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12391__A0 cpu.DM0.readdata\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07937__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11162_ net2561 net160 net414 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
XANTENNA__10941__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__C net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__and2_1
X_11093_ cpu.RF0.registers\[2\]\[23\] net152 net422 vssd1 vssd1 vccd1 vccd1 _00527_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12143__B1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ cpu.IM0.address_IM\[17\] _05306_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__nor2_1
XANTENNA__08898__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 _01501_ vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11185__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13230__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08362__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 cpu.f0.write_data\[30\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 cpu.LCD0.lcd_rs vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 cpu.f0.write_data\[11\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net88 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ clknet_leaf_90_clk _00916_ net1276 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11995_ net505 _05766_ _05912_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_55_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11913__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ clknet_leaf_4_clk _00847_ net1150 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10946_ net1556 net927 _05685_ net275 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_clk_X clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13380__CLK clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13665_ clknet_leaf_63_clk _00778_ net1308 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ cpu.DM0.readdata\[14\] _05086_ net737 vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12948__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12749__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ net2291 cpu.LCD0.row_2\[10\] net999 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
XANTENNA__09075__A0 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13596_ clknet_leaf_8_clk _00709_ net1165 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _01869_ _01873_ _01889_ _06311_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a31o_1
XANTENNA__10224__A3 _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_67_clk_X clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12478_ _01798_ _06268_ _06269_ net263 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09378__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ clknet_leaf_105_clk _01330_ net1155 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11429_ net2018 net149 net383 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10117__X _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__B1 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_96_clk _01261_ net1231 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10932__A1 _04517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06970_ cpu.RF0.registers\[16\]\[25\] net582 net573 cpu.RF0.registers\[9\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a22o_1
X_14079_ clknet_leaf_106_clk _01192_ net1140 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12134__B1 _06034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09354__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_2
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_1
X_08640_ cpu.IM0.address_IM\[3\] net554 _03929_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_
+ sky130_fd_sc_hd__a22o_2
XANTENNA__09550__B2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1092 net1094 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XANTENNA__10160__A2 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ cpu.RF0.registers\[8\]\[5\] _02014_ net658 cpu.RF0.registers\[13\]\[5\] _03849_
+ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_46_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11823__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08105__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07522_ net1058 cpu.RF0.registers\[22\]\[6\] net802 vssd1 vssd1 vccd1 vccd1 _02813_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload89_A clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ cpu.RF0.registers\[16\]\[1\] net582 _02728_ _02730_ _02735_ vssd1 vssd1 vccd1
+ vccd1 _02744_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_100_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06404_ cpu.f0.i\[30\] vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07384_ cpu.RF0.registers\[13\]\[2\] net598 _02648_ _02657_ _02665_ vssd1 vssd1 vccd1
+ vccd1 _02675_ sky130_fd_sc_hd__a2111o_1
X_09123_ net302 _04381_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07040__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout317_A _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ net1028 cpu.RF0.registers\[31\]\[31\] net825 vssd1 vssd1 vccd1 vccd1 _04345_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13103__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07092__A2 _02381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14229__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ cpu.RF0.registers\[16\]\[28\] net635 _03274_ _03275_ _03281_ vssd1 vssd1
+ vccd1 vccd1 _03296_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09369__A1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold520 cpu.RF0.registers\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09248__B net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold531 cpu.RF0.registers\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 cpu.RF0.registers\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12373__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 cpu.RF0.registers\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 cpu.RF0.registers\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 cpu.RF0.registers\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 cpu.RF0.registers\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 cpu.RF0.registers\[31\]\[0\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14379__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _05235_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or2_1
XANTENNA__12125__B1 _06025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06888__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ _04196_ _04197_ net439 vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a21oi_2
X_09887_ _05173_ _05174_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or2_1
Xhold1220 cpu.RF0.registers\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 cpu.RF0.registers\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net1075 cpu.RF0.registers\[17\]\[16\] net882 vssd1 vssd1 vccd1 vccd1 _04129_
+ sky130_fd_sc_hd__and3_1
Xhold1242 cpu.RF0.registers\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 cpu.RF0.registers\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 cpu.RF0.registers\[4\]\[16\] vssd1 vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 cpu.RF0.registers\[21\]\[4\] vssd1 vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1286 cpu.RF0.registers\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1297 cpu.RF0.registers\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ net1095 cpu.RF0.registers\[24\]\[18\] net871 vssd1 vssd1 vccd1 vccd1 _04060_
+ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_37_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ net993 _04663_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ net2110 net175 net340 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07304__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07512__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ net987 cpu.f0.data_adr\[5\] vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13450_ clknet_leaf_102_clk _00563_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ cpu.LCD0.row_1\[68\] cpu.LCD0.row_1\[76\] net904 vssd1 vssd1 vccd1 vccd1
+ _00292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12401_ cpu.DM0.data_i\[9\] net515 _06222_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a21o_1
XANTENNA__07607__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12600__A1 cpu.SR1.char_in\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ clknet_leaf_9_clk _00494_ net1163 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ _05685_ cpu.LCD0.row_1\[7\] net896 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ cpu.LCD0.cnt_20ms\[9\] cpu.LCD0.cnt_20ms\[8\] _06202_ cpu.LCD0.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07083__A2 _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ cpu.LCD0.row_1\[14\] _05994_ _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ clknet_leaf_70_clk _01115_ net1326 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11214_ net2222 net201 net407 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
X_12194_ cpu.LCD0.row_2\[91\] _05983_ _06011_ cpu.LCD0.row_2\[51\] vssd1 vssd1 vccd1
+ vccd1 _06092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__11908__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_11145_ net2673 net222 net416 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__09780__B2 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__12116__B1 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_94_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ cpu.RF0.registers\[2\]\[6\] net231 net423 vssd1 vssd1 vccd1 vccd1 _00510_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13746__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08335__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _05289_ _05302_ _05300_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10142__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A cpu.IM0.address_IM\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07125__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11643__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__B _03233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ net1730 net174 net316 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__mux2_1
XANTENNA__08518__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_74_clk _00830_ net1324 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10929_ cpu.DM0.readdata\[29\] _04551_ net738 vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13126__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_75_clk _00761_ net1321 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13579_ clknet_leaf_90_clk _00692_ net1279 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07795__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08253__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_47_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13276__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14521__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12206__C _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08540__X _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 net309 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XANTENNA__11818__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ net449 _04509_ _04692_ _02758_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__o211a_1
XANTENNA__08574__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 _05941_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_6
Xfanout329 _05939_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_6
XANTENNA__12107__B1 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _04027_ _04028_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a21oi_1
X_06953_ cpu.RF0.registers\[20\]\[26\] net594 _02226_ _02231_ net621 vssd1 vssd1 vccd1
+ vccd1 _02244_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06501__A cpu.K0.keyvalid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _02830_ _03833_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__xor2_1
XANTENNA__07316__B _02606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ net966 net801 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__and2_4
XANTENNA__10133__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ net950 cpu.RF0.registers\[14\]\[3\] net840 vssd1 vssd1 vccd1 vccd1 _03914_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07035__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11553__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ net1107 cpu.RF0.registers\[31\]\[5\] net858 vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07505_ net306 _02794_ _02760_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__or3b_1
XANTENNA__07332__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ net1106 cpu.RF0.registers\[25\]\[7\] net864 vssd1 vssd1 vccd1 vccd1 _03776_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ net976 cpu.RF0.registers\[10\]\[1\] net789 vssd1 vssd1 vccd1 vccd1 _02727_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_80_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14051__CLK clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07367_ net976 cpu.RF0.registers\[11\]\[2\] net777 vssd1 vssd1 vccd1 vccd1 _02658_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout601_A _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12594__A0 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13619__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1343_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _04391_ _04395_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_21_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08163__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ cpu.RF0.registers\[10\]\[4\] net570 net566 cpu.RF0.registers\[11\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09037_ net952 cpu.RF0.registers\[15\]\[31\] net825 vssd1 vssd1 vccd1 vccd1 _04328_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09211__A0 _03402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 _01674_ vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 a1.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13769__CLK clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout970_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 cpu.RF0.registers\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 cpu.SR1.char_in\[7\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 cpu.RF0.registers\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10372__A2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout830 _02129_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
Xfanout841 _02049_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_70_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout852 _02038_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_6
X_09939_ cpu.IM0.address_IM\[8\] net933 _05222_ _05223_ vssd1 vssd1 vccd1 vccd1 _00031_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_70_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_8
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
XANTENNA__09514__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14401__Q cpu.IG0.Instr\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout896 net901 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_4
X_12950_ clknet_leaf_20_clk _00139_ net1168 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1050 _01633_ vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ net2594 net243 net323 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
Xhold1061 cpu.RF0.registers\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09722__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__A_N cpu.IM0.address_IM\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1072 cpu.RF0.registers\[6\]\[0\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 _00311_ vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_1_clk cpu.c0.next_count\[12\] net1137 vssd1 vssd1 vccd1 vccd1
+ cpu.c0.count\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 cpu.LCD0.cnt_500hz\[7\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11463__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14620_ clknet_leaf_30_clk _01721_ net1209 vssd1 vssd1 vccd1 vccd1 cpu.f0.write_data\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11832_ net2036 net253 net333 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__mux2_1
XANTENNA__09278__A0 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13149__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14551_ clknet_leaf_56_clk net2127 net1370 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11763_ net2408 net131 net342 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10832__A0 cpu.DM0.readdata\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10714_ a1.BUSY_O cpu.RU0.state\[2\] net929 _00016_ vssd1 vssd1 vccd1 vccd1 _05686_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ clknet_leaf_83_clk _00615_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14482_ clknet_leaf_30_clk net1410 net1209 vssd1 vssd1 vccd1 vccd1 cpu.RU0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ net1969 net144 net353 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13433_ clknet_leaf_91_clk _00546_ net1277 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13299__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ net2407 net2431 net900 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
XANTENNA__14544__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A0 _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ clknet_leaf_70_clk _00477_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10576_ _05675_ cpu.LCD0.row_1\[0\] net896 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
X_12315_ net1369 _05946_ _06196_ _05957_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__a31o_1
XANTENNA__10060__A1 cpu.IM0.address_IM\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13295_ clknet_leaf_33_clk cpu.RU0.next_FetchedData\[2\] net1248 vssd1 vssd1 vccd1
+ vccd1 cpu.DM0.data_i\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12246_ cpu.LCD0.row_2\[37\] _06004_ _06006_ cpu.LCD0.row_1\[37\] _06141_ vssd1 vssd1
+ vccd1 vccd1 _06142_ sky130_fd_sc_hd__a221o_1
XANTENNA__08801__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11638__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07213__C1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ cpu.LCD0.nextState\[1\] net743 net557 _06007_ cpu.LCD0.row_2\[114\] vssd1
+ vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11128_ net2355 net160 net418 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09505__A1 _03629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ net2100 _05827_ net426 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09632__A _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08248__A _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14074__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10823__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ cpu.RF0.registers\[5\]\[15\] net703 _03559_ _03560_ vssd1 vssd1 vccd1 vccd1
+ _03561_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07295__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07221_ net1035 cpu.RF0.registers\[24\]\[9\] net811 vssd1 vssd1 vccd1 vccd1 _02512_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07047__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ net1044 cpu.RF0.registers\[21\]\[11\] net798 vssd1 vssd1 vccd1 vccd1 _02443_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08414__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13911__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09992__A1 cpu.IM0.address_IM\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07083_ cpu.RF0.registers\[5\]\[18\] _02148_ _02354_ _02358_ _02367_ vssd1 vssd1
+ vccd1 vccd1 _02374_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_93_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11548__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08547__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11000__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06558__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__C_N _04601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 _05148_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_2
Xfanout148 net151 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
Xfanout159 _05832_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_07985_ net1094 cpu.RF0.registers\[31\]\[28\] net857 vssd1 vssd1 vccd1 vccd1 _03276_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04808_ _05009_ _05014_ net277 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a2bb2o_1
X_06936_ net1029 cpu.RF0.registers\[18\]\[26\] net769 vssd1 vssd1 vccd1 vccd1 _02227_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _02436_ net300 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__xor2_1
XANTENNA__14417__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ net962 cpu.RF0.registers\[7\]\[27\] net817 vssd1 vssd1 vccd1 vccd1 _02158_
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__B1 cpu.IM0.address_IM\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _03886_ _03888_ _03893_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__or4_1
X_09586_ _04384_ _04781_ _04872_ net486 _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_06798_ cpu.IM0.address_IM\[30\] net551 _02088_ _02081_ vssd1 vssd1 vccd1 vccd1 _02089_
+ sky130_fd_sc_hd__a22o_2
XANTENNA__07062__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ cpu.RF0.registers\[31\]\[6\] net686 net670 cpu.RF0.registers\[22\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a22o_1
XANTENNA__10975__X _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout816_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A0 cpu.f0.data_adr\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13441__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08468_ net951 cpu.RF0.registers\[15\]\[8\] net857 vssd1 vssd1 vccd1 vccd1 _03759_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07286__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ cpu.RF0.registers\[18\]\[0\] net579 _02707_ _02708_ _02709_ vssd1 vssd1 vccd1
+ vccd1 _02710_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ cpu.RF0.registers\[3\]\[10\] net643 _03671_ _03672_ _03681_ vssd1 vssd1 vccd1
+ vccd1 _03690_ sky130_fd_sc_hd__a2111o_1
X_10430_ cpu.f0.i\[27\] net268 vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13591__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10042__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09983__A1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__B cpu.IG0.Instr\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ cpu.f0.i\[27\] _05582_ cpu.f0.i\[28\] vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13300__Q cpu.DM0.data_i\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06797__A1 cpu.RF0.registers\[0\]\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ _05984_ net743 _05996_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ clknet_leaf_48_clk _00260_ net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[44\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_72_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10292_ _05534_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_72_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08538__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11458__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net2861 _05945_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
Xhold180 cpu.f0.write_data\[14\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 cpu.RF0.registers\[26\]\[13\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12815__RESET_B net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__B1 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 _02053_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_89_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout671 _02045_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_89_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12098__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout682 net683 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13982_ clknet_leaf_84_clk _01095_ net1270 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout693 _02026_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_6
X_12933_ clknet_leaf_29_clk _00122_ net1201 vssd1 vssd1 vccd1 vccd1 a1.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11193__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12864_ clknet_leaf_16_clk _00083_ net1196 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14603_ clknet_leaf_54_clk net2345 net1349 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_11815_ net1725 net191 net334 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ net2573 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10805__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14534_ clknet_leaf_45_clk _01636_ net1311 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[45\]
+ sky130_fd_sc_hd__dfstp_1
X_11746_ net2313 net193 net343 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__mux2_1
XANTENNA__12270__A2 _06006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13934__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07700__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14465_ clknet_leaf_22_clk _01575_ net1174 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_11677_ net1650 net201 net351 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ net2358 net2283 net897 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
X_13416_ clknet_leaf_85_clk _00529_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14396_ clknet_leaf_21_clk _01507_ net1176 vssd1 vssd1 vccd1 vccd1 cpu.IG0.Instr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10033__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ clknet_leaf_79_clk _00460_ net1316 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[0\]\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_10559_ net56 net920 vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10584__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A _03145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13278_ clknet_leaf_19_clk cpu.RU0.next_FetchedInstr\[17\] net1176 vssd1 vssd1 vccd1
+ vccd1 cpu.FetchedInstr\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08529__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12229_ cpu.LCD0.row_2\[68\] _05988_ _05998_ cpu.LCD0.row_2\[12\] vssd1 vssd1 vccd1
+ vccd1 _06126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07737__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13314__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07770_ cpu.RF0.registers\[4\]\[21\] net586 net582 cpu.RF0.registers\[16\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a22o_1
XANTENNA__06986__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06721_ net1081 cpu.RF0.registers\[20\]\[30\] net874 vssd1 vssd1 vccd1 vccd1 _02012_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09440_ _04497_ _04724_ _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__o21bai_2
XANTENNA__08701__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06652_ net1422 net892 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[20\] sky130_fd_sc_hd__and2_1
XANTENNA__09081__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09371_ _04415_ _04655_ _04661_ _04653_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__o211a_1
XANTENNA__10795__X _05744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06583_ cpu.LCD0.cnt_500hz\[11\] _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__nand2_1
XANTENNA__11831__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ net1086 cpu.RF0.registers\[25\]\[12\] net862 vssd1 vssd1 vccd1 vccd1 _03613_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_99_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12261__A2 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload71_A clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08253_ net1092 cpu.RF0.registers\[17\]\[15\] net884 vssd1 vssd1 vccd1 vccd1 _03544_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07204_ cpu.RF0.registers\[8\]\[10\] net611 _02476_ _02477_ _02479_ vssd1 vssd1 vccd1
+ vccd1 _02495_ sky130_fd_sc_hd__a2111o_1
XANTENNA_wire774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08184_ net444 _03472_ _03473_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__nand3_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07135_ cpu.RF0.registers\[21\]\[15\] net593 _02425_ net623 vssd1 vssd1 vccd1 vccd1
+ _02426_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1041_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07976__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ net974 cpu.RF0.registers\[3\]\[18\] net823 vssd1 vssd1 vccd1 vccd1 _02357_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08441__A _03729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1306_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12182__D1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09824__X _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14132__RESET_B net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ cpu.RF0.registers\[25\]\[29\] net648 _03241_ _03248_ _03249_ vssd1 vssd1
+ vccd1 vccd1 _03259_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06896__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ net450 _03992_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nor2_1
X_06919_ net742 _02208_ cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout933_A _01787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07899_ cpu.RF0.registers\[15\]\[29\] _02167_ _03189_ net623 vssd1 vssd1 vccd1 vccd1
+ _03190_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09638_ _02384_ net441 vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13957__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__C net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _04594_ _04711_ _04750_ net480 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07223__C net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net2534 net238 net361 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XANTENNA__11741__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12580_ cpu.DM0.data_i\[4\] _06339_ cpu.DM0.data_i\[5\] vssd1 vssd1 vccd1 vccd1 _06343_
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__12252__A2 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10865__B _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08616__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11531_ net1793 net137 net370 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__mux2_1
XANTENNA__10802__A3 _05748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12981__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ clknet_leaf_100_clk _01363_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11462_ net1591 net148 net381 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XANTENNA__09405__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08903__X _04194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ clknet_leaf_70_clk _00381_ net1329 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10413_ net1124 _05624_ net264 net1978 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08054__C _02062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ clknet_leaf_9_clk _01294_ net1166 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11393_ net1903 net180 net387 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__mux2_1
X_13132_ clknet_leaf_50_clk net2680 net1383 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_10344_ _05578_ _05579_ net308 vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__or3b_1
XANTENNA__13337__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11188__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13063_ clknet_leaf_47_clk _00243_ net1354 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09166__B _03766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ cpu.f0.i\[15\] _05518_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12014_ net2151 net186 net312 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10105__B cpu.IM0.address_IM\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_2
XFILLER_0_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13965_ clknet_leaf_101_clk _01078_ net1212 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08144__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ clknet_leaf_25_clk _00105_ net1186 vssd1 vssd1 vccd1 vccd1 cpu.f0.num\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload8_A clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_98_clk _01009_ net1269 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ clknet_leaf_31_clk _00066_ net1204 vssd1 vssd1 vccd1 vccd1 cpu.f0.data_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11651__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__A2 _06022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ net2909 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ clknet_leaf_49_clk _01619_ net1359 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_2\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11729_ net1911 net136 net346 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ clknet_leaf_27_clk _01558_ net1187 vssd1 vssd1 vccd1 vccd1 cpu.f0.i\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09947__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14379_ clknet_leaf_33_clk _01490_ net1247 vssd1 vssd1 vccd1 vccd1 cpu.CU0.opcode\[6\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold905 cpu.LCD0.row_1\[98\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 cpu.RF0.registers\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 cpu.LCD0.row_1\[55\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 cpu.LCD0.row_2\[114\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 cpu.RF0.registers\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11098__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ _04228_ _04229_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09791__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ _04160_ _04161_ _04159_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ cpu.RF0.registers\[28\]\[22\] net578 _03093_ _03103_ _03104_ vssd1 vssd1
+ vccd1 vccd1 _03113_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11826__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ net523 _03041_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__o21ai_4
X_06704_ _01949_ _01944_ cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_write_i
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07684_ cpu.RF0.registers\[26\]\[16\] net599 _02952_ _02959_ _02961_ vssd1 vssd1
+ vccd1 vccd1 _02975_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _04414_ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and2_1
X_06635_ a1.CPU_DAT_O\[3\] net895 vssd1 vssd1 vccd1 vccd1 cpu.RU0.next_FetchedInstr\[3\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07043__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11561__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ net298 _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__nand2_1
X_06566_ _01944_ _01946_ _01949_ cpu.RU0.state\[0\] vssd1 vssd1 vccd1 vccd1 _01950_
+ sky130_fd_sc_hd__or4b_1
XANTENNA__08438__A1 cpu.IM0.address_IM\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ _02832_ _02868_ _02903_ net490 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a31o_1
XANTENNA__10245__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09285_ _04574_ _04575_ _04565_ _04568_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__a211o_1
X_06497_ cpu.DM0.dhit cpu.f0.state\[7\] _01887_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a21o_1
XANTENNA__07110__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10796__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ _03522_ _03524_ _03526_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14605__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12392__S net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ net1099 cpu.RF0.registers\[20\]\[20\] net875 vssd1 vssd1 vccd1 vccd1 _03458_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07118_ net545 _02385_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__or2_1
XANTENNA__09267__A _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ cpu.RF0.registers\[28\]\[22\] net705 net684 cpu.RF0.registers\[24\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout883_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ cpu.RF0.registers\[17\]\[19\] net605 _02317_ _02320_ _02323_ vssd1 vssd1
+ vccd1 vccd1 _02340_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1309_X net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ cpu.IM0.address_IM\[18\] net932 _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _00041_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09273__Y _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _02470_ net516 _05852_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21o_1
X_13750_ clknet_leaf_71_clk _00863_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12701_ net1897 net2199 net1004 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ clknet_leaf_79_clk _00794_ net1321 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10893_ net1670 net188 net431 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
XANTENNA__14135__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12632_ cpu.LCD0.row_2\[34\] net1584 net999 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__mux2_1
XANTENNA__12225__A2 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08346__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _01874_ _06314_ _06322_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or4_4
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11984__A1 _05822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14302_ clknet_leaf_83_clk _01415_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11514_ net1970 net200 net370 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__mux2_1
X_12494_ cpu.f0.i\[14\] _06277_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nand2_1
XANTENNA__14285__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ clknet_leaf_14_clk _01346_ net1256 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11445_ net2802 net214 net379 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11736__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ clknet_leaf_71_clk _01277_ net1338 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11376_ net1910 net224 net387 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__mux2_1
XANTENNA__08081__A _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13115_ clknet_leaf_46_clk net2601 net1360 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_10327_ _05479_ _05563_ _05565_ net724 cpu.f0.data_adr\[24\] vssd1 vssd1 vccd1 vccd1
+ _00077_ sky130_fd_sc_hd__o32a_1
X_14095_ clknet_leaf_83_clk _01208_ net1275 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13046_ clknet_leaf_54_clk _00226_ net1352 vssd1 vssd1 vccd1 vccd1 cpu.LCD0.row_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10258_ _01805_ _05500_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and2_1
XANTENNA__12877__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1230 net1232 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11646__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1241 net1268 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1252 net1254 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_4
X_10189_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__or2_1
Xfanout1263 net1265 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1274 net1275 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1285 net1287 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1296 net1299 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__clkbuf_2
X_13948_ clknet_leaf_15_clk _01061_ net1244 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10786__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ clknet_leaf_65_clk _00992_ net1282 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11381__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06420_ _01777_ _01830_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12216__A2 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07798__C net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__A1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07160__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14628__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10778__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12209__C _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09070_ _03195_ _03197_ _03233_ net488 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07643__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ net1097 cpu.RF0.registers\[17\]\[24\] net884 vssd1 vssd1 vccd1 vccd1 _03312_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13652__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 cpu.RF0.registers\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold713 cpu.RF0.registers\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 cpu.LCD0.row_1\[9\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold735 cpu.LCD0.row_2\[71\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 a1.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 cpu.RF0.registers\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__C net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold768 _01616_ vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ cpu.IM0.address_IM\[11\] _05242_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__and2_1
Xhold779 cpu.LCD0.row_1\[46\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08923_ net938 cpu.RF0.registers\[7\]\[27\] net844 vssd1 vssd1 vccd1 vccd1 _04214_
+ sky130_fd_sc_hd__and3_1
XANTENNA__07038__C net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__Y _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1402 cpu.RF0.registers\[1\]\[10\] vssd1 vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ _04132_ _04136_ _04140_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or4_1
Xhold1413 cpu.RF0.registers\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1004_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1424 cpu.RF0.registers\[0\]\[0\] vssd1 vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06877__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1435 cpu.LCD0.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 cpu.RF0.registers\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net2852 sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ net1031 cpu.RF0.registers\[19\]\[22\] net820 vssd1 vssd1 vccd1 vccd1 _03096_
+ sky130_fd_sc_hd__and3_1
Xhold1457 cpu.RF0.registers\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ cpu.RF0.registers\[29\]\[18\] net673 net667 _04063_ _04066_ vssd1 vssd1 vccd1
+ vccd1 _04076_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_93_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1468 cpu.RF0.registers\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net2874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1479 cpu.RF0.registers\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net2885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14158__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ cpu.RF0.registers\[18\]\[20\] net579 net574 cpu.RF0.registers\[9\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__a22o_1
X_07667_ net1024 cpu.RF0.registers\[23\]\[16\] net816 vssd1 vssd1 vccd1 vccd1 _02958_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11291__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__B net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ _04401_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06618_ _01977_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nor2_1
XANTENNA__08166__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ net968 cpu.RF0.registers\[14\]\[12\] net762 vssd1 vssd1 vccd1 vccd1 _02889_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10218__A1 cpu.f0.data_adr\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07070__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__B2 cpu.f0.i\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06549_ _01780_ net1129 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__nand2_1
X_09337_ _04619_ _04622_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07095__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ net445 net291 _02311_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ net443 _03507_ _03508_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09199_ _04482_ _04489_ _04479_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21o_1
XANTENNA__12416__A cpu.DM0.data_i\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net2391 net151 net407 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XANTENNA__09387__A2 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14404__Q cpu.IG0.Instr\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ net1960 net177 net415 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10941__A2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ cpu.IM0.address_IM\[23\] _02310_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__nand2_1
X_11092_ net2165 net164 net422 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XANTENNA__11466__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10043_ cpu.IM0.address_IM\[17\] _05306_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__and2_1
Xhold40 cpu.LCD0.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 cpu.FetchedInstr\[14\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 cpu.FetchedInstr\[19\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 net93 vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 cpu.f0.data_adr\[11\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _00175_ vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13802_ clknet_leaf_100_clk _00915_ net1217 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11994_ net1754 net128 net314 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13525__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_103_clk _00846_ net1214 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10945_ net1683 net926 _05683_ net274 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ clknet_leaf_3_clk _00777_ net1160 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ net1855 net200 net430 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
X_12615_ net2416 net2376 net1007 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XANTENNA__07411__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09075__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13595_ clknet_leaf_12_clk _00708_ net1226 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12546_ _06312_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__nor2_1
XANTENNA__14235__RESET_B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _01798_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__nand2_1
XANTENNA_4 _05753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_99_clk _01329_ net1233 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11428_ net1596 net156 net382 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__B2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14147_ clknet_leaf_77_clk _01260_ net1318 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11359_ cpu.RF0.registers\[10\]\[23\] net153 net390 vssd1 vssd1 vccd1 vccd1 _00783_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10393__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14078_ clknet_leaf_85_clk _01191_ net1271 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13055__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ clknet_leaf_54_clk _00001_ vssd1 vssd1 vccd1 vccd1 cpu.LCD0.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_2
Xfanout1071 cpu.IG0.Instr\[21\] vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_6_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1091 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_2
Xfanout1093 net1094 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
X_08570_ cpu.RF0.registers\[21\]\[5\] net647 net641 cpu.RF0.registers\[19\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06994__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07521_ net1056 cpu.RF0.registers\[23\]\[6\] net818 vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__and3_1
XANTENNA__10448__B2 a1.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14450__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ net978 cpu.RF0.registers\[6\]\[1\] net803 vssd1 vssd1 vccd1 vccd1 _02743_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12000__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07864__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06403_ net2916 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07383_ cpu.RF0.registers\[28\]\[2\] net577 _02653_ _02661_ _02663_ vssd1 vssd1 vccd1
+ vccd1 _02674_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09066__A1 cpu.RF0.registers\[0\]\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__C net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ net484 _04409_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__X _03564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ net1027 cpu.RF0.registers\[26\]\[31\] net786 vssd1 vssd1 vccd1 vccd1 _04344_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload100_A clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ cpu.RF0.registers\[25\]\[28\] _02059_ net640 cpu.RF0.registers\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold510 cpu.RF0.registers\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10867__A1_N net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold521 cpu.c0.count\[2\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold532 cpu.RF0.registers\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13958__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold543 cpu.RF0.registers\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold554 cpu.RF0.registers\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08041__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 cpu.RF0.registers\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09816__Y _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_A cpu.DM0.ihit vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold576 cpu.RF0.registers\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 cpu.RF0.registers\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 cpu.RF0.registers\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _05214_ _05215_ _05226_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__o31a_2
XANTENNA__07991__C net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11286__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06888__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A _02037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net490 _04195_ _03019_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10136__B1 cpu.IM0.address_IM\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _05173_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__nand2_1
Xhold1210 cpu.DM0.readdata\[25\] vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 cpu.f0.state\[0\] vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07065__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 cpu.RF0.registers\[17\]\[20\] vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ _04090_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nand2_1
Xhold1243 cpu.RF0.registers\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 cpu.LCD0.row_1\[91\] vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1265 cpu.c0.count\[6\] vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 cpu.RF0.registers\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 a1.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 cpu.RF0.registers\[14\]\[1\] vssd1 vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ net1100 cpu.RF0.registers\[22\]\[18\] _02038_ vssd1 vssd1 vccd1 vccd1 _04059_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ cpu.RF0.registers\[12\]\[17\] net572 _02996_ _03001_ _03006_ vssd1 vssd1
+ vccd1 vccd1 _03010_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_0_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _03976_ _03977_ _03984_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__or4_4
XANTENNA__13698__CLK clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10730_ net993 _05073_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ net2253 cpu.LCD0.row_1\[75\] net898 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11034__B cpu.IG0.Instr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ net2712 net733 _06223_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__o21a_1
X_13380_ clknet_leaf_100_clk _00493_ net1229 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ net995 _02579_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10873__B _04774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12331_ net1446 _06203_ _06205_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ net745 _05987_ _05993_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3_1
XANTENNA__13078__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__C net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14001_ clknet_leaf_77_clk _01114_ net1332 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08568__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ net2580 net212 net407 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12193_ cpu.LCD0.row_2\[35\] _06004_ _06028_ cpu.LCD0.row_1\[115\] _06090_ vssd1
+ vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__a221o_1
XANTENNA__14323__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__09455__A _02982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net1818 net224 net415 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XANTENNA__12116__A1 cpu.LCD0.row_1\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12116__B2 cpu.LCD0.row_2\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__11196__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06594__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09174__B _03899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11075_ cpu.RF0.registers\[2\]\[5\] net233 net423 vssd1 vssd1 vccd1 vccd1 _00509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _05289_ _05300_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__or3_1
XANTENNA__14473__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__C net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ net2378 net195 net316 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13716_ clknet_leaf_71_clk _00829_ net1330 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07846__A2 _02160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928_ net1649 net146 net432 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13647_ clknet_leaf_86_clk _00760_ net1274 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10859_ _05229_ _05789_ net720 vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09189__X _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13578_ clknet_leaf_100_clk _00691_ net1216 vssd1 vssd1 vccd1 vccd1 cpu.RF0.registers\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12529_ cpu.f0.i\[28\] _06299_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13369__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_2
Xfanout319 _05941_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
X_09740_ _04027_ _04028_ net494 vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__o21ai_1
X_06952_ _02239_ _02240_ _02241_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__or4_1
.ends

