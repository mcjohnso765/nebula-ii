VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO team_04
  CLASS BLOCK ;
  FOREIGN team_04 ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 500.000 ;
  PIN ACK_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 466.990 496.000 467.270 500.000 ;
    END
  END ACK_I
  PIN ADR_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 518.510 496.000 518.790 500.000 ;
    END
  END ADR_O[0]
  PIN ADR_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 212.610 496.000 212.890 500.000 ;
    END
  END ADR_O[10]
  PIN ADR_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 496.000 216.110 500.000 ;
    END
  END ADR_O[11]
  PIN ADR_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END ADR_O[12]
  PIN ADR_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 444.450 496.000 444.730 500.000 ;
    END
  END ADR_O[13]
  PIN ADR_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 183.630 496.000 183.910 500.000 ;
    END
  END ADR_O[14]
  PIN ADR_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.190 496.000 177.470 500.000 ;
    END
  END ADR_O[15]
  PIN ADR_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 460.550 496.000 460.830 500.000 ;
    END
  END ADR_O[16]
  PIN ADR_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 450.890 496.000 451.170 500.000 ;
    END
  END ADR_O[17]
  PIN ADR_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 515.290 496.000 515.570 500.000 ;
    END
  END ADR_O[18]
  PIN ADR_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 496.000 135.610 500.000 ;
    END
  END ADR_O[19]
  PIN ADR_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 370.390 496.000 370.670 500.000 ;
    END
  END ADR_O[1]
  PIN ADR_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 496.000 122.730 500.000 ;
    END
  END ADR_O[20]
  PIN ADR_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 496.000 80.870 500.000 ;
    END
  END ADR_O[21]
  PIN ADR_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 496.000 71.210 500.000 ;
    END
  END ADR_O[22]
  PIN ADR_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 496.000 42.230 500.000 ;
    END
  END ADR_O[23]
  PIN ADR_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 331.750 496.000 332.030 500.000 ;
    END
  END ADR_O[24]
  PIN ADR_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 260.910 496.000 261.190 500.000 ;
    END
  END ADR_O[25]
  PIN ADR_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 280.230 496.000 280.510 500.000 ;
    END
  END ADR_O[26]
  PIN ADR_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 286.670 496.000 286.950 500.000 ;
    END
  END ADR_O[27]
  PIN ADR_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 312.430 496.000 312.710 500.000 ;
    END
  END ADR_O[28]
  PIN ADR_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 328.530 496.000 328.810 500.000 ;
    END
  END ADR_O[29]
  PIN ADR_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 351.070 496.000 351.350 500.000 ;
    END
  END ADR_O[2]
  PIN ADR_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 373.610 496.000 373.890 500.000 ;
    END
  END ADR_O[30]
  PIN ADR_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 309.210 496.000 309.490 500.000 ;
    END
  END ADR_O[31]
  PIN ADR_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 383.270 496.000 383.550 500.000 ;
    END
  END ADR_O[3]
  PIN ADR_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END ADR_O[4]
  PIN ADR_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 325.310 496.000 325.590 500.000 ;
    END
  END ADR_O[5]
  PIN ADR_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 302.770 496.000 303.050 500.000 ;
    END
  END ADR_O[6]
  PIN ADR_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 496.000 299.830 500.000 ;
    END
  END ADR_O[7]
  PIN ADR_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 244.810 496.000 245.090 500.000 ;
    END
  END ADR_O[8]
  PIN ADR_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 267.350 496.000 267.630 500.000 ;
    END
  END ADR_O[9]
  PIN CYC_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 496.000 167.810 500.000 ;
    END
  END CYC_O
  PIN DAT_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 438.010 496.000 438.290 500.000 ;
    END
  END DAT_I[0]
  PIN DAT_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 316.240 550.000 316.840 ;
    END
  END DAT_I[10]
  PIN DAT_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 363.840 550.000 364.440 ;
    END
  END DAT_I[11]
  PIN DAT_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 380.840 550.000 381.440 ;
    END
  END DAT_I[12]
  PIN DAT_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 431.570 496.000 431.850 500.000 ;
    END
  END DAT_I[13]
  PIN DAT_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 374.040 550.000 374.640 ;
    END
  END DAT_I[14]
  PIN DAT_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 391.040 550.000 391.640 ;
    END
  END DAT_I[15]
  PIN DAT_I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 353.640 550.000 354.240 ;
    END
  END DAT_I[16]
  PIN DAT_I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 319.640 550.000 320.240 ;
    END
  END DAT_I[17]
  PIN DAT_I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 326.440 550.000 327.040 ;
    END
  END DAT_I[18]
  PIN DAT_I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 329.840 550.000 330.440 ;
    END
  END DAT_I[19]
  PIN DAT_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 412.250 496.000 412.530 500.000 ;
    END
  END DAT_I[1]
  PIN DAT_I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 350.240 550.000 350.840 ;
    END
  END DAT_I[20]
  PIN DAT_I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 336.640 550.000 337.240 ;
    END
  END DAT_I[21]
  PIN DAT_I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 346.840 550.000 347.440 ;
    END
  END DAT_I[22]
  PIN DAT_I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 425.130 496.000 425.410 500.000 ;
    END
  END DAT_I[23]
  PIN DAT_I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 323.040 550.000 323.640 ;
    END
  END DAT_I[24]
  PIN DAT_I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 401.240 550.000 401.840 ;
    END
  END DAT_I[25]
  PIN DAT_I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 340.040 550.000 340.640 ;
    END
  END DAT_I[26]
  PIN DAT_I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 377.440 550.000 378.040 ;
    END
  END DAT_I[27]
  PIN DAT_I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 434.790 496.000 435.070 500.000 ;
    END
  END DAT_I[28]
  PIN DAT_I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 367.240 550.000 367.840 ;
    END
  END DAT_I[29]
  PIN DAT_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 428.350 496.000 428.630 500.000 ;
    END
  END DAT_I[2]
  PIN DAT_I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 360.440 550.000 361.040 ;
    END
  END DAT_I[30]
  PIN DAT_I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 357.040 550.000 357.640 ;
    END
  END DAT_I[31]
  PIN DAT_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 418.690 496.000 418.970 500.000 ;
    END
  END DAT_I[3]
  PIN DAT_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 408.040 550.000 408.640 ;
    END
  END DAT_I[4]
  PIN DAT_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 404.640 550.000 405.240 ;
    END
  END DAT_I[5]
  PIN DAT_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 415.470 496.000 415.750 500.000 ;
    END
  END DAT_I[6]
  PIN DAT_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 421.910 496.000 422.190 500.000 ;
    END
  END DAT_I[7]
  PIN DAT_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 333.240 550.000 333.840 ;
    END
  END DAT_I[8]
  PIN DAT_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 343.440 550.000 344.040 ;
    END
  END DAT_I[9]
  PIN DAT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 231.240 550.000 231.840 ;
    END
  END DAT_O[0]
  PIN DAT_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 312.840 550.000 313.440 ;
    END
  END DAT_O[10]
  PIN DAT_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END DAT_O[11]
  PIN DAT_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END DAT_O[12]
  PIN DAT_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END DAT_O[13]
  PIN DAT_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END DAT_O[14]
  PIN DAT_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END DAT_O[15]
  PIN DAT_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 272.040 550.000 272.640 ;
    END
  END DAT_O[16]
  PIN DAT_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END DAT_O[17]
  PIN DAT_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END DAT_O[18]
  PIN DAT_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END DAT_O[19]
  PIN DAT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END DAT_O[1]
  PIN DAT_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 238.040 550.000 238.640 ;
    END
  END DAT_O[20]
  PIN DAT_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 261.840 550.000 262.440 ;
    END
  END DAT_O[21]
  PIN DAT_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END DAT_O[22]
  PIN DAT_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END DAT_O[23]
  PIN DAT_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 241.440 550.000 242.040 ;
    END
  END DAT_O[24]
  PIN DAT_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 268.640 550.000 269.240 ;
    END
  END DAT_O[25]
  PIN DAT_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 258.440 550.000 259.040 ;
    END
  END DAT_O[26]
  PIN DAT_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 255.040 550.000 255.640 ;
    END
  END DAT_O[27]
  PIN DAT_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 244.840 550.000 245.440 ;
    END
  END DAT_O[28]
  PIN DAT_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 248.240 550.000 248.840 ;
    END
  END DAT_O[29]
  PIN DAT_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END DAT_O[2]
  PIN DAT_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END DAT_O[30]
  PIN DAT_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END DAT_O[31]
  PIN DAT_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END DAT_O[3]
  PIN DAT_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END DAT_O[4]
  PIN DAT_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END DAT_O[5]
  PIN DAT_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END DAT_O[6]
  PIN DAT_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END DAT_O[7]
  PIN DAT_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END DAT_O[8]
  PIN DAT_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END DAT_O[9]
  PIN SEL_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 367.170 496.000 367.450 500.000 ;
    END
  END SEL_O[0]
  PIN SEL_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 380.050 496.000 380.330 500.000 ;
    END
  END SEL_O[1]
  PIN SEL_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 389.710 496.000 389.990 500.000 ;
    END
  END SEL_O[2]
  PIN SEL_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END SEL_O[3]
  PIN STB_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 496.000 164.590 500.000 ;
    END
  END STB_O
  PIN WE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 399.370 496.000 399.650 500.000 ;
    END
  END WE_O
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 392.930 496.000 393.210 500.000 ;
    END
  END en
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END gpio_in[33]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.190 496.000 16.470 500.000 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END gpio_in[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 409.030 496.000 409.310 500.000 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 496.000 232.210 500.000 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 454.110 496.000 454.390 500.000 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 496.000 39.010 500.000 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 496.000 61.550 500.000 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 496.000 32.570 500.000 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 496.000 74.430 500.000 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 496.000 171.030 500.000 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 496.000 154.930 500.000 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 496.000 58.330 500.000 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 496.000 22.910 500.000 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 496.000 10.030 500.000 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 496.000 64.770 500.000 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 496.000 129.170 500.000 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 496.000 193.570 500.000 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 496.000 35.790 500.000 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 496.000 77.650 500.000 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 496.000 235.430 500.000 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 496.000 45.450 500.000 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 495.970 496.000 496.250 500.000 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 496.000 180.690 500.000 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 499.190 496.000 499.470 500.000 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 470.210 496.000 470.490 500.000 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 496.000 84.090 500.000 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 457.330 496.000 457.610 500.000 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 531.390 496.000 531.670 500.000 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 521.730 496.000 522.010 500.000 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 496.000 145.270 500.000 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 496.000 19.690 500.000 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 431.840 550.000 432.440 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 496.000 187.130 500.000 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 496.000 0.370 500.000 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 524.950 496.000 525.230 500.000 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 496.000 251.530 500.000 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 512.070 496.000 512.350 500.000 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 270.570 496.000 270.850 500.000 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 496.000 6.810 500.000 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 496.000 48.670 500.000 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 496.000 87.310 500.000 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 496.000 3.590 500.000 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 496.000 151.710 500.000 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 496.000 238.650 500.000 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 496.000 158.150 500.000 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 496.000 125.950 500.000 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 496.000 116.290 500.000 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 447.670 496.000 447.950 500.000 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 402.590 496.000 402.870 500.000 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 544.270 496.000 544.550 500.000 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 496.000 174.250 500.000 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 405.810 496.000 406.090 500.000 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 496.000 90.530 500.000 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 496.000 132.390 500.000 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 496.000 248.310 500.000 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 496.000 225.770 500.000 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 496.000 26.130 500.000 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 496.000 103.410 500.000 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 463.770 496.000 464.050 500.000 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 496.000 29.350 500.000 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 500.000 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 496.000 148.490 500.000 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 496.000 51.890 500.000 ;
    END
  END gpio_out[33]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 357.510 496.000 357.790 500.000 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 496.000 161.370 500.000 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 496.000 13.250 500.000 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 496.000 93.750 500.000 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 496.000 67.990 500.000 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 496.000 55.110 500.000 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 496.000 142.050 500.000 ;
    END
  END gpio_out[9]
  PIN mem_adr_start[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 360.730 496.000 361.010 500.000 ;
    END
  END mem_adr_start[0]
  PIN mem_adr_start[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 441.230 496.000 441.510 500.000 ;
    END
  END mem_adr_start[10]
  PIN mem_adr_start[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 222.270 496.000 222.550 500.000 ;
    END
  END mem_adr_start[11]
  PIN mem_adr_start[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 199.730 496.000 200.010 500.000 ;
    END
  END mem_adr_start[12]
  PIN mem_adr_start[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 190.070 496.000 190.350 500.000 ;
    END
  END mem_adr_start[13]
  PIN mem_adr_start[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 500.000 ;
    END
  END mem_adr_start[14]
  PIN mem_adr_start[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 534.610 496.000 534.890 500.000 ;
    END
  END mem_adr_start[15]
  PIN mem_adr_start[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 489.530 496.000 489.810 500.000 ;
    END
  END mem_adr_start[16]
  PIN mem_adr_start[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 508.850 496.000 509.130 500.000 ;
    END
  END mem_adr_start[17]
  PIN mem_adr_start[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 547.490 496.000 547.770 500.000 ;
    END
  END mem_adr_start[18]
  PIN mem_adr_start[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.550 496.000 138.830 500.000 ;
    END
  END mem_adr_start[19]
  PIN mem_adr_start[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 363.950 496.000 364.230 500.000 ;
    END
  END mem_adr_start[1]
  PIN mem_adr_start[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 505.630 496.000 505.910 500.000 ;
    END
  END mem_adr_start[20]
  PIN mem_adr_start[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 486.310 496.000 486.590 500.000 ;
    END
  END mem_adr_start[21]
  PIN mem_adr_start[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 502.410 496.000 502.690 500.000 ;
    END
  END mem_adr_start[22]
  PIN mem_adr_start[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 528.170 496.000 528.450 500.000 ;
    END
  END mem_adr_start[23]
  PIN mem_adr_start[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 254.470 496.000 254.750 500.000 ;
    END
  END mem_adr_start[24]
  PIN mem_adr_start[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 257.690 496.000 257.970 500.000 ;
    END
  END mem_adr_start[25]
  PIN mem_adr_start[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 277.010 496.000 277.290 500.000 ;
    END
  END mem_adr_start[26]
  PIN mem_adr_start[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 273.790 496.000 274.070 500.000 ;
    END
  END mem_adr_start[27]
  PIN mem_adr_start[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 305.990 496.000 306.270 500.000 ;
    END
  END mem_adr_start[28]
  PIN mem_adr_start[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 315.650 496.000 315.930 500.000 ;
    END
  END mem_adr_start[29]
  PIN mem_adr_start[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 344.630 496.000 344.910 500.000 ;
    END
  END mem_adr_start[2]
  PIN mem_adr_start[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 496.000 296.610 500.000 ;
    END
  END mem_adr_start[30]
  PIN mem_adr_start[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 293.110 496.000 293.390 500.000 ;
    END
  END mem_adr_start[31]
  PIN mem_adr_start[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 496.000 338.470 500.000 ;
    END
  END mem_adr_start[3]
  PIN mem_adr_start[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 322.090 496.000 322.370 500.000 ;
    END
  END mem_adr_start[4]
  PIN mem_adr_start[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 318.870 496.000 319.150 500.000 ;
    END
  END mem_adr_start[5]
  PIN mem_adr_start[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 289.890 496.000 290.170 500.000 ;
    END
  END mem_adr_start[6]
  PIN mem_adr_start[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.450 496.000 283.730 500.000 ;
    END
  END mem_adr_start[7]
  PIN mem_adr_start[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 241.590 496.000 241.870 500.000 ;
    END
  END mem_adr_start[8]
  PIN mem_adr_start[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.130 496.000 264.410 500.000 ;
    END
  END mem_adr_start[9]
  PIN memory_size[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 476.650 496.000 476.930 500.000 ;
    END
  END memory_size[0]
  PIN memory_size[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 396.150 496.000 396.430 500.000 ;
    END
  END memory_size[10]
  PIN memory_size[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 219.050 496.000 219.330 500.000 ;
    END
  END memory_size[11]
  PIN memory_size[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.390 496.000 209.670 500.000 ;
    END
  END memory_size[12]
  PIN memory_size[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 496.000 206.450 500.000 ;
    END
  END memory_size[13]
  PIN memory_size[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 541.050 496.000 541.330 500.000 ;
    END
  END memory_size[14]
  PIN memory_size[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 473.430 496.000 473.710 500.000 ;
    END
  END memory_size[15]
  PIN memory_size[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 119.230 496.000 119.510 500.000 ;
    END
  END memory_size[16]
  PIN memory_size[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.790 496.000 113.070 500.000 ;
    END
  END memory_size[17]
  PIN memory_size[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.350 496.000 106.630 500.000 ;
    END
  END memory_size[18]
  PIN memory_size[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 96.690 496.000 96.970 500.000 ;
    END
  END memory_size[19]
  PIN memory_size[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 354.290 496.000 354.570 500.000 ;
    END
  END memory_size[1]
  PIN memory_size[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 496.000 109.850 500.000 ;
    END
  END memory_size[20]
  PIN memory_size[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.910 496.000 100.190 500.000 ;
    END
  END memory_size[21]
  PIN memory_size[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 537.830 496.000 538.110 500.000 ;
    END
  END memory_size[22]
  PIN memory_size[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 479.870 496.000 480.150 500.000 ;
    END
  END memory_size[23]
  PIN memory_size[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 483.090 496.000 483.370 500.000 ;
    END
  END memory_size[24]
  PIN memory_size[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 492.750 496.000 493.030 500.000 ;
    END
  END memory_size[25]
  PIN memory_size[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 386.490 496.000 386.770 500.000 ;
    END
  END memory_size[26]
  PIN memory_size[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.970 496.000 335.250 500.000 ;
    END
  END memory_size[27]
  PIN memory_size[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 347.850 496.000 348.130 500.000 ;
    END
  END memory_size[28]
  PIN memory_size[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END memory_size[29]
  PIN memory_size[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 435.240 550.000 435.840 ;
    END
  END memory_size[2]
  PIN memory_size[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END memory_size[30]
  PIN memory_size[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END memory_size[31]
  PIN memory_size[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 438.640 550.000 439.240 ;
    END
  END memory_size[3]
  PIN memory_size[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 442.040 550.000 442.640 ;
    END
  END memory_size[4]
  PIN memory_size[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 445.440 550.000 446.040 ;
    END
  END memory_size[5]
  PIN memory_size[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END memory_size[6]
  PIN memory_size[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END memory_size[7]
  PIN memory_size[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END memory_size[8]
  PIN memory_size[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END memory_size[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 546.000 27.240 550.000 27.840 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 487.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 544.370 487.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 486.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 547.790 489.220 ;
      LAYER met2 ;
        RECT 0.650 495.720 3.030 496.810 ;
        RECT 3.870 495.720 6.250 496.810 ;
        RECT 7.090 495.720 9.470 496.810 ;
        RECT 10.310 495.720 12.690 496.810 ;
        RECT 13.530 495.720 15.910 496.810 ;
        RECT 16.750 495.720 19.130 496.810 ;
        RECT 19.970 495.720 22.350 496.810 ;
        RECT 23.190 495.720 25.570 496.810 ;
        RECT 26.410 495.720 28.790 496.810 ;
        RECT 29.630 495.720 32.010 496.810 ;
        RECT 32.850 495.720 35.230 496.810 ;
        RECT 36.070 495.720 38.450 496.810 ;
        RECT 39.290 495.720 41.670 496.810 ;
        RECT 42.510 495.720 44.890 496.810 ;
        RECT 45.730 495.720 48.110 496.810 ;
        RECT 48.950 495.720 51.330 496.810 ;
        RECT 52.170 495.720 54.550 496.810 ;
        RECT 55.390 495.720 57.770 496.810 ;
        RECT 58.610 495.720 60.990 496.810 ;
        RECT 61.830 495.720 64.210 496.810 ;
        RECT 65.050 495.720 67.430 496.810 ;
        RECT 68.270 495.720 70.650 496.810 ;
        RECT 71.490 495.720 73.870 496.810 ;
        RECT 74.710 495.720 77.090 496.810 ;
        RECT 77.930 495.720 80.310 496.810 ;
        RECT 81.150 495.720 83.530 496.810 ;
        RECT 84.370 495.720 86.750 496.810 ;
        RECT 87.590 495.720 89.970 496.810 ;
        RECT 90.810 495.720 93.190 496.810 ;
        RECT 94.030 495.720 96.410 496.810 ;
        RECT 97.250 495.720 99.630 496.810 ;
        RECT 100.470 495.720 102.850 496.810 ;
        RECT 103.690 495.720 106.070 496.810 ;
        RECT 106.910 495.720 109.290 496.810 ;
        RECT 110.130 495.720 112.510 496.810 ;
        RECT 113.350 495.720 115.730 496.810 ;
        RECT 116.570 495.720 118.950 496.810 ;
        RECT 119.790 495.720 122.170 496.810 ;
        RECT 123.010 495.720 125.390 496.810 ;
        RECT 126.230 495.720 128.610 496.810 ;
        RECT 129.450 495.720 131.830 496.810 ;
        RECT 132.670 495.720 135.050 496.810 ;
        RECT 135.890 495.720 138.270 496.810 ;
        RECT 139.110 495.720 141.490 496.810 ;
        RECT 142.330 495.720 144.710 496.810 ;
        RECT 145.550 495.720 147.930 496.810 ;
        RECT 148.770 495.720 151.150 496.810 ;
        RECT 151.990 495.720 154.370 496.810 ;
        RECT 155.210 495.720 157.590 496.810 ;
        RECT 158.430 495.720 160.810 496.810 ;
        RECT 161.650 495.720 164.030 496.810 ;
        RECT 164.870 495.720 167.250 496.810 ;
        RECT 168.090 495.720 170.470 496.810 ;
        RECT 171.310 495.720 173.690 496.810 ;
        RECT 174.530 495.720 176.910 496.810 ;
        RECT 177.750 495.720 180.130 496.810 ;
        RECT 180.970 495.720 183.350 496.810 ;
        RECT 184.190 495.720 186.570 496.810 ;
        RECT 187.410 495.720 189.790 496.810 ;
        RECT 190.630 495.720 193.010 496.810 ;
        RECT 193.850 495.720 196.230 496.810 ;
        RECT 197.070 495.720 199.450 496.810 ;
        RECT 200.290 495.720 202.670 496.810 ;
        RECT 203.510 495.720 205.890 496.810 ;
        RECT 206.730 495.720 209.110 496.810 ;
        RECT 209.950 495.720 212.330 496.810 ;
        RECT 213.170 495.720 215.550 496.810 ;
        RECT 216.390 495.720 218.770 496.810 ;
        RECT 219.610 495.720 221.990 496.810 ;
        RECT 222.830 495.720 225.210 496.810 ;
        RECT 226.050 495.720 228.430 496.810 ;
        RECT 229.270 495.720 231.650 496.810 ;
        RECT 232.490 495.720 234.870 496.810 ;
        RECT 235.710 495.720 238.090 496.810 ;
        RECT 238.930 495.720 241.310 496.810 ;
        RECT 242.150 495.720 244.530 496.810 ;
        RECT 245.370 495.720 247.750 496.810 ;
        RECT 248.590 495.720 250.970 496.810 ;
        RECT 251.810 495.720 254.190 496.810 ;
        RECT 255.030 495.720 257.410 496.810 ;
        RECT 258.250 495.720 260.630 496.810 ;
        RECT 261.470 495.720 263.850 496.810 ;
        RECT 264.690 495.720 267.070 496.810 ;
        RECT 267.910 495.720 270.290 496.810 ;
        RECT 271.130 495.720 273.510 496.810 ;
        RECT 274.350 495.720 276.730 496.810 ;
        RECT 277.570 495.720 279.950 496.810 ;
        RECT 280.790 495.720 283.170 496.810 ;
        RECT 284.010 495.720 286.390 496.810 ;
        RECT 287.230 495.720 289.610 496.810 ;
        RECT 290.450 495.720 292.830 496.810 ;
        RECT 293.670 495.720 296.050 496.810 ;
        RECT 296.890 495.720 299.270 496.810 ;
        RECT 300.110 495.720 302.490 496.810 ;
        RECT 303.330 495.720 305.710 496.810 ;
        RECT 306.550 495.720 308.930 496.810 ;
        RECT 309.770 495.720 312.150 496.810 ;
        RECT 312.990 495.720 315.370 496.810 ;
        RECT 316.210 495.720 318.590 496.810 ;
        RECT 319.430 495.720 321.810 496.810 ;
        RECT 322.650 495.720 325.030 496.810 ;
        RECT 325.870 495.720 328.250 496.810 ;
        RECT 329.090 495.720 331.470 496.810 ;
        RECT 332.310 495.720 334.690 496.810 ;
        RECT 335.530 495.720 337.910 496.810 ;
        RECT 338.750 495.720 341.130 496.810 ;
        RECT 341.970 495.720 344.350 496.810 ;
        RECT 345.190 495.720 347.570 496.810 ;
        RECT 348.410 495.720 350.790 496.810 ;
        RECT 351.630 495.720 354.010 496.810 ;
        RECT 354.850 495.720 357.230 496.810 ;
        RECT 358.070 495.720 360.450 496.810 ;
        RECT 361.290 495.720 363.670 496.810 ;
        RECT 364.510 495.720 366.890 496.810 ;
        RECT 367.730 495.720 370.110 496.810 ;
        RECT 370.950 495.720 373.330 496.810 ;
        RECT 374.170 495.720 376.550 496.810 ;
        RECT 377.390 495.720 379.770 496.810 ;
        RECT 380.610 495.720 382.990 496.810 ;
        RECT 383.830 495.720 386.210 496.810 ;
        RECT 387.050 495.720 389.430 496.810 ;
        RECT 390.270 495.720 392.650 496.810 ;
        RECT 393.490 495.720 395.870 496.810 ;
        RECT 396.710 495.720 399.090 496.810 ;
        RECT 399.930 495.720 402.310 496.810 ;
        RECT 403.150 495.720 405.530 496.810 ;
        RECT 406.370 495.720 408.750 496.810 ;
        RECT 409.590 495.720 411.970 496.810 ;
        RECT 412.810 495.720 415.190 496.810 ;
        RECT 416.030 495.720 418.410 496.810 ;
        RECT 419.250 495.720 421.630 496.810 ;
        RECT 422.470 495.720 424.850 496.810 ;
        RECT 425.690 495.720 428.070 496.810 ;
        RECT 428.910 495.720 431.290 496.810 ;
        RECT 432.130 495.720 434.510 496.810 ;
        RECT 435.350 495.720 437.730 496.810 ;
        RECT 438.570 495.720 440.950 496.810 ;
        RECT 441.790 495.720 444.170 496.810 ;
        RECT 445.010 495.720 447.390 496.810 ;
        RECT 448.230 495.720 450.610 496.810 ;
        RECT 451.450 495.720 453.830 496.810 ;
        RECT 454.670 495.720 457.050 496.810 ;
        RECT 457.890 495.720 460.270 496.810 ;
        RECT 461.110 495.720 463.490 496.810 ;
        RECT 464.330 495.720 466.710 496.810 ;
        RECT 467.550 495.720 469.930 496.810 ;
        RECT 470.770 495.720 473.150 496.810 ;
        RECT 473.990 495.720 476.370 496.810 ;
        RECT 477.210 495.720 479.590 496.810 ;
        RECT 480.430 495.720 482.810 496.810 ;
        RECT 483.650 495.720 486.030 496.810 ;
        RECT 486.870 495.720 489.250 496.810 ;
        RECT 490.090 495.720 492.470 496.810 ;
        RECT 493.310 495.720 495.690 496.810 ;
        RECT 496.530 495.720 498.910 496.810 ;
        RECT 499.750 495.720 502.130 496.810 ;
        RECT 502.970 495.720 505.350 496.810 ;
        RECT 506.190 495.720 508.570 496.810 ;
        RECT 509.410 495.720 511.790 496.810 ;
        RECT 512.630 495.720 515.010 496.810 ;
        RECT 515.850 495.720 518.230 496.810 ;
        RECT 519.070 495.720 521.450 496.810 ;
        RECT 522.290 495.720 524.670 496.810 ;
        RECT 525.510 495.720 527.890 496.810 ;
        RECT 528.730 495.720 531.110 496.810 ;
        RECT 531.950 495.720 534.330 496.810 ;
        RECT 535.170 495.720 537.550 496.810 ;
        RECT 538.390 495.720 540.770 496.810 ;
        RECT 541.610 495.720 543.990 496.810 ;
        RECT 544.830 495.720 547.210 496.810 ;
        RECT 0.100 4.280 547.760 495.720 ;
        RECT 0.650 4.000 3.030 4.280 ;
        RECT 3.870 4.000 6.250 4.280 ;
        RECT 7.090 4.000 9.470 4.280 ;
        RECT 10.310 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.970 4.280 ;
        RECT 90.810 4.000 93.190 4.280 ;
        RECT 94.030 4.000 96.410 4.280 ;
        RECT 97.250 4.000 99.630 4.280 ;
        RECT 100.470 4.000 102.850 4.280 ;
        RECT 103.690 4.000 202.670 4.280 ;
        RECT 203.510 4.000 221.990 4.280 ;
        RECT 222.830 4.000 254.190 4.280 ;
        RECT 255.030 4.000 263.850 4.280 ;
        RECT 264.690 4.000 267.070 4.280 ;
        RECT 267.910 4.000 276.730 4.280 ;
        RECT 277.570 4.000 279.950 4.280 ;
        RECT 280.790 4.000 312.150 4.280 ;
        RECT 312.990 4.000 325.030 4.280 ;
        RECT 325.870 4.000 334.690 4.280 ;
        RECT 335.530 4.000 547.760 4.280 ;
      LAYER met3 ;
        RECT 3.990 480.440 546.000 487.045 ;
        RECT 4.400 479.040 546.000 480.440 ;
        RECT 3.990 453.240 546.000 479.040 ;
        RECT 4.400 451.840 546.000 453.240 ;
        RECT 3.990 446.440 546.000 451.840 ;
        RECT 3.990 445.040 545.600 446.440 ;
        RECT 3.990 443.040 546.000 445.040 ;
        RECT 3.990 441.640 545.600 443.040 ;
        RECT 3.990 439.640 546.000 441.640 ;
        RECT 3.990 438.240 545.600 439.640 ;
        RECT 3.990 436.240 546.000 438.240 ;
        RECT 4.400 434.840 545.600 436.240 ;
        RECT 3.990 432.840 546.000 434.840 ;
        RECT 4.400 431.440 545.600 432.840 ;
        RECT 3.990 429.440 546.000 431.440 ;
        RECT 4.400 428.040 546.000 429.440 ;
        RECT 3.990 409.040 546.000 428.040 ;
        RECT 3.990 407.640 545.600 409.040 ;
        RECT 3.990 405.640 546.000 407.640 ;
        RECT 3.990 404.240 545.600 405.640 ;
        RECT 3.990 402.240 546.000 404.240 ;
        RECT 3.990 400.840 545.600 402.240 ;
        RECT 3.990 392.040 546.000 400.840 ;
        RECT 3.990 390.640 545.600 392.040 ;
        RECT 3.990 381.840 546.000 390.640 ;
        RECT 3.990 380.440 545.600 381.840 ;
        RECT 3.990 378.440 546.000 380.440 ;
        RECT 3.990 377.040 545.600 378.440 ;
        RECT 3.990 375.040 546.000 377.040 ;
        RECT 3.990 373.640 545.600 375.040 ;
        RECT 3.990 368.240 546.000 373.640 ;
        RECT 3.990 366.840 545.600 368.240 ;
        RECT 3.990 364.840 546.000 366.840 ;
        RECT 3.990 363.440 545.600 364.840 ;
        RECT 3.990 361.440 546.000 363.440 ;
        RECT 3.990 360.040 545.600 361.440 ;
        RECT 3.990 358.040 546.000 360.040 ;
        RECT 3.990 356.640 545.600 358.040 ;
        RECT 3.990 354.640 546.000 356.640 ;
        RECT 3.990 353.240 545.600 354.640 ;
        RECT 3.990 351.240 546.000 353.240 ;
        RECT 3.990 349.840 545.600 351.240 ;
        RECT 3.990 347.840 546.000 349.840 ;
        RECT 3.990 346.440 545.600 347.840 ;
        RECT 3.990 344.440 546.000 346.440 ;
        RECT 3.990 343.040 545.600 344.440 ;
        RECT 3.990 341.040 546.000 343.040 ;
        RECT 3.990 339.640 545.600 341.040 ;
        RECT 3.990 337.640 546.000 339.640 ;
        RECT 3.990 336.240 545.600 337.640 ;
        RECT 3.990 334.240 546.000 336.240 ;
        RECT 3.990 332.840 545.600 334.240 ;
        RECT 3.990 330.840 546.000 332.840 ;
        RECT 3.990 329.440 545.600 330.840 ;
        RECT 3.990 327.440 546.000 329.440 ;
        RECT 3.990 326.040 545.600 327.440 ;
        RECT 3.990 324.040 546.000 326.040 ;
        RECT 3.990 322.640 545.600 324.040 ;
        RECT 3.990 320.640 546.000 322.640 ;
        RECT 3.990 319.240 545.600 320.640 ;
        RECT 3.990 317.240 546.000 319.240 ;
        RECT 3.990 315.840 545.600 317.240 ;
        RECT 3.990 313.840 546.000 315.840 ;
        RECT 3.990 312.440 545.600 313.840 ;
        RECT 3.990 310.440 546.000 312.440 ;
        RECT 4.400 309.040 546.000 310.440 ;
        RECT 3.990 296.840 546.000 309.040 ;
        RECT 4.400 295.440 546.000 296.840 ;
        RECT 3.990 273.040 546.000 295.440 ;
        RECT 3.990 271.640 545.600 273.040 ;
        RECT 3.990 269.640 546.000 271.640 ;
        RECT 4.400 268.240 545.600 269.640 ;
        RECT 3.990 262.840 546.000 268.240 ;
        RECT 3.990 261.440 545.600 262.840 ;
        RECT 3.990 259.440 546.000 261.440 ;
        RECT 3.990 258.040 545.600 259.440 ;
        RECT 3.990 256.040 546.000 258.040 ;
        RECT 4.400 254.640 545.600 256.040 ;
        RECT 3.990 249.240 546.000 254.640 ;
        RECT 3.990 247.840 545.600 249.240 ;
        RECT 3.990 245.840 546.000 247.840 ;
        RECT 4.400 244.440 545.600 245.840 ;
        RECT 3.990 242.440 546.000 244.440 ;
        RECT 4.400 241.040 545.600 242.440 ;
        RECT 3.990 239.040 546.000 241.040 ;
        RECT 4.400 237.640 545.600 239.040 ;
        RECT 3.990 235.640 546.000 237.640 ;
        RECT 4.400 234.240 546.000 235.640 ;
        RECT 3.990 232.240 546.000 234.240 ;
        RECT 4.400 230.840 545.600 232.240 ;
        RECT 3.990 228.840 546.000 230.840 ;
        RECT 4.400 227.440 546.000 228.840 ;
        RECT 3.990 225.440 546.000 227.440 ;
        RECT 4.400 224.040 546.000 225.440 ;
        RECT 3.990 222.040 546.000 224.040 ;
        RECT 4.400 220.640 546.000 222.040 ;
        RECT 3.990 218.640 546.000 220.640 ;
        RECT 4.400 217.240 546.000 218.640 ;
        RECT 3.990 198.240 546.000 217.240 ;
        RECT 4.400 196.840 546.000 198.240 ;
        RECT 3.990 28.240 546.000 196.840 ;
        RECT 3.990 26.840 545.600 28.240 ;
        RECT 3.990 10.715 546.000 26.840 ;
      LAYER met4 ;
        RECT 23.295 12.415 23.940 458.825 ;
        RECT 26.340 12.415 174.240 458.825 ;
        RECT 176.640 12.415 177.540 458.825 ;
        RECT 179.940 12.415 327.840 458.825 ;
        RECT 330.240 12.415 331.140 458.825 ;
        RECT 333.540 12.415 481.440 458.825 ;
        RECT 483.840 12.415 484.740 458.825 ;
        RECT 487.140 12.415 519.505 458.825 ;
  END
END team_04
END LIBRARY

