* NGSPICE file created from team_02_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt team_02_Wrapper gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36] gpio_in[37] gpio_in[3] gpio_in[4]
+ gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10]
+ gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17]
+ gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23]
+ gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2]
+ gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34] gpio_oeb[35] gpio_oeb[36]
+ gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8]
+ gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14]
+ gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20]
+ gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27]
+ gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33]
+ gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3] gpio_out[4] gpio_out[5]
+ gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1] irq[2] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1
+ wb_clk_i wb_rst_i wbm_ack_i wbm_adr_o[0] wbm_adr_o[10] wbm_adr_o[11] wbm_adr_o[12]
+ wbm_adr_o[13] wbm_adr_o[14] wbm_adr_o[15] wbm_adr_o[16] wbm_adr_o[17] wbm_adr_o[18]
+ wbm_adr_o[19] wbm_adr_o[1] wbm_adr_o[20] wbm_adr_o[21] wbm_adr_o[22] wbm_adr_o[23]
+ wbm_adr_o[24] wbm_adr_o[25] wbm_adr_o[26] wbm_adr_o[27] wbm_adr_o[28] wbm_adr_o[29]
+ wbm_adr_o[2] wbm_adr_o[30] wbm_adr_o[31] wbm_adr_o[3] wbm_adr_o[4] wbm_adr_o[5]
+ wbm_adr_o[6] wbm_adr_o[7] wbm_adr_o[8] wbm_adr_o[9] wbm_cyc_o wbm_dat_i[0] wbm_dat_i[10]
+ wbm_dat_i[11] wbm_dat_i[12] wbm_dat_i[13] wbm_dat_i[14] wbm_dat_i[15] wbm_dat_i[16]
+ wbm_dat_i[17] wbm_dat_i[18] wbm_dat_i[19] wbm_dat_i[1] wbm_dat_i[20] wbm_dat_i[21]
+ wbm_dat_i[22] wbm_dat_i[23] wbm_dat_i[24] wbm_dat_i[25] wbm_dat_i[26] wbm_dat_i[27]
+ wbm_dat_i[28] wbm_dat_i[29] wbm_dat_i[2] wbm_dat_i[30] wbm_dat_i[31] wbm_dat_i[3]
+ wbm_dat_i[4] wbm_dat_i[5] wbm_dat_i[6] wbm_dat_i[7] wbm_dat_i[8] wbm_dat_i[9] wbm_dat_o[0]
+ wbm_dat_o[10] wbm_dat_o[11] wbm_dat_o[12] wbm_dat_o[13] wbm_dat_o[14] wbm_dat_o[15]
+ wbm_dat_o[16] wbm_dat_o[17] wbm_dat_o[18] wbm_dat_o[19] wbm_dat_o[1] wbm_dat_o[20]
+ wbm_dat_o[21] wbm_dat_o[22] wbm_dat_o[23] wbm_dat_o[24] wbm_dat_o[25] wbm_dat_o[26]
+ wbm_dat_o[27] wbm_dat_o[28] wbm_dat_o[29] wbm_dat_o[2] wbm_dat_o[30] wbm_dat_o[31]
+ wbm_dat_o[3] wbm_dat_o[4] wbm_dat_o[5] wbm_dat_o[6] wbm_dat_o[7] wbm_dat_o[8] wbm_dat_o[9]
+ wbm_sel_o[0] wbm_sel_o[1] wbm_sel_o[2] wbm_sel_o[3] wbm_stb_o wbm_we_o wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_103_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09671_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] net869 net865 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08731__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ net973 _04381_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08553_ net101 net1660 net893 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XANTENNA__13083__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818__1372 vssd1 vssd1 vccd1 vccd1 _16818__1372/HI net1372 sky130_fd_sc_hd__conb_1
XANTENNA__08428__B net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07504_ net1648 team_02_WB.instance_to_wrap.ramload\[1\] net968 vssd1 vssd1 vccd1
+ vccd1 _02830_ sky130_fd_sc_hd__mux2_1
X_08484_ _04311_ _04312_ net742 net751 net1732 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1071_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1169_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09105_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] net725 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a221o_1
XANTENNA__08798__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16746__1300 vssd1 vssd1 vccd1 vccd1 _16746__1300/HI net1300 sky130_fd_sc_hd__conb_1
X_09036_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] net721 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\]
+ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold340 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 team_02_WB.instance_to_wrap.top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 net1760
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12897__A2 _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold373 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09762__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold395 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout820 _04650_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_8
XANTENNA__15741__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\] net815 net803 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a22o_1
Xfanout842 _04672_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout853 _04655_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_8
Xfanout864 _04647_ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_4
Xfanout875 _04668_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09514__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 _04632_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
X_09869_ _05526_ _05528_ _05530_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__or4_2
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
Xhold1040 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11744__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1062 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net233 net1791 net546 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1073 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
X_16702__1256 vssd1 vssd1 vccd1 vccd1 _16702__1256/HI net1256 sky130_fd_sc_hd__conb_1
X_12880_ team_02_WB.instance_to_wrap.top.pc\[9\] _05635_ vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1084 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15891__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ net353 net2224 net552 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14550_ net1105 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
X_11762_ net347 net2563 net561 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03353_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ _06356_ _06363_ net391 vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13374__B1_N _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ net1028 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XANTENNA__12575__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ net335 net2651 net568 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
X_16220_ clknet_leaf_37_wb_clk_i _02665_ _01177_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13260__A _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input92_A wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\] _03300_ vssd1 vssd1 vccd1
+ vccd1 _03314_ sky130_fd_sc_hd__nor2_1
X_10644_ team_02_WB.instance_to_wrap.top.pc\[19\] _06255_ _06295_ vssd1 vssd1 vccd1
+ vccd1 _06296_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16151_ clknet_leaf_38_wb_clk_i net1626 _01109_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10575_ team_02_WB.instance_to_wrap.top.pc\[29\] _06225_ vssd1 vssd1 vccd1 vccd1
+ _06227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ team_02_WB.instance_to_wrap.top.a1.row1\[107\] _03216_ _03240_ team_02_WB.instance_to_wrap.top.a1.row2\[11\]
+ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__a221o_1
XANTENNA__10596__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15102_ clknet_leaf_4_wb_clk_i _01553_ _00060_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15271__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ net304 net2670 net503 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
XANTENNA__10060__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16082_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[0\] _01040_
+ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__dfrtp_1
X_13294_ _03178_ _03184_ _03195_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o211ai_1
XANTENNA_output179_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ net1169 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12245_ net281 net2176 net510 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09185__A _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12176_ net276 net2158 net517 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11127_ net403 _06529_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09505__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ net441 _06676_ _06677_ net428 _06692_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[22\]
+ sky130_fd_sc_hd__a221o_1
X_15935_ clknet_leaf_29_wb_clk_i _02386_ _00893_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_60_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11654__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] net732 net672 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a22o_1
X_15866_ clknet_leaf_120_wb_clk_i _02317_ _00824_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14817_ net1203 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15797_ clknet_leaf_124_wb_clk_i _02248_ _00755_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13065__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14748_ net1182 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12485__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ net1167 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16418_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[17\]
+ _01292_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire597_A _05790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15614__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ clknet_leaf_101_wb_clk_i _02782_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10051__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11829__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15764__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11000__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07984_ _03872_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__or2_1
XANTENNA__11839__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] net823 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12500__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout377_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09654_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] net656 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _04386_ _04400_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15144__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ _05249_ _05251_ _05253_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__or4_4
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08536_ net88 net1622 net892 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08873__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12395__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ team_02_WB.instance_to_wrap.top.a1.data\[0\] net916 vssd1 vssd1 vccd1 vccd1
+ _04320_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout711_A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15294__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10290__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14904__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10360_ _05793_ _06012_ _05749_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09983__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _04701_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__or2_2
XFILLER_0_104_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10291_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] net789 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a221o_1
X_12030_ net347 net1801 net469 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XANTENNA__09196__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13239__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[15\] vssd1 vssd1 vccd1
+ vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_02_WB.START_ADDR_VAL_REG\[5\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold192 net146 vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16641__1212 vssd1 vssd1 vccd1 vccd1 _16641__1212/HI net1212 sky130_fd_sc_hd__conb_1
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_8
Xfanout661 _04480_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
Xfanout672 _04475_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_8
Xfanout683 _04471_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_2
X_13981_ net1030 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
Xfanout694 _04467_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_6
XANTENNA__11474__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15720_ clknet_leaf_57_wb_clk_i _02171_ _00678_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12932_ _02886_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__and2_1
XANTENNA__08349__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15651_ clknet_leaf_40_wb_clk_i _02102_ _00609_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ _03402_ _06254_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__nand2_1
X_14602_ net1178 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
X_11814_ net303 net2292 net554 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15582_ clknet_leaf_4_wb_clk_i _02033_ _00540_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11058__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ _07408_ _07417_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__nor2_1
XANTENNA__15637__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09120__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14533_ net1089 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11745_ net281 net2093 net560 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ net1072 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
X_11676_ net277 net2706 net570 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ clknet_leaf_30_wb_clk_i _02648_ _01160_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13415_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _03300_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10627_ team_02_WB.instance_to_wrap.top.pc\[14\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _06279_ sky130_fd_sc_hd__or2_1
X_14395_ net1060 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14814__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10033__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16134_ clknet_leaf_7_wb_clk_i net1550 _01092_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09908__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13346_ team_02_WB.instance_to_wrap.top.a1.row1\[1\] _03227_ _03238_ team_02_WB.instance_to_wrap.top.a1.row2\[33\]
+ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10558_ _04826_ _06210_ _06141_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11649__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ clknet_leaf_1_wb_clk_i _02516_ _01023_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ _03178_ _03188_ _03174_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10489_ _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15016_ net1168 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16817__1371 vssd1 vssd1 vccd1 vccd1 _16817__1371/HI net1371 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12228_ net340 net2253 net514 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
XANTENNA__09726__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ net331 net2642 net521 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16412__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15918_ clknet_leaf_40_wb_clk_i _02369_ _00876_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ clknet_leaf_29_wb_clk_i _02300_ _00807_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09370_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] net734 net728 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\]
+ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16562__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ _04194_ _04196_ _04188_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08252_ _04131_ _04132_ _04106_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__or3b_4
XFILLER_0_6_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08183_ _04053_ net224 _04050_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13210__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10024__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__A _05461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701__1255 vssd1 vssd1 vccd1 vccd1 _16701__1255/HI net1255 sky130_fd_sc_hd__conb_1
XFILLER_0_3_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput220 net220 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09178__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13059__B net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07967_ _03841_ _03850_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a21o_2
XANTENNA__10699__A _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout759_A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\] net658 net633 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\]
+ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07898_ _03772_ _03782_ _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a21oi_2
X_09637_ _05301_ _05302_ _05304_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout926_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09568_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] net702 net675 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08519_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09499_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] net735 net650 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a22o_1
XANTENNA__08616__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07520__B net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ _06002_ _06006_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ net408 _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ team_02_WB.START_ADDR_VAL_REG\[8\] _04356_ vssd1 vssd1 vccd1 vccd1 net222
+ sky130_fd_sc_hd__and2_1
X_10412_ _05012_ net367 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nand2_1
X_11392_ _06095_ _06097_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__nand2_1
XANTENNA__09956__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ net1143 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XANTENNA__08632__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13131_ _00005_ team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[4\] sky130_fd_sc_hd__or2_1
X_10343_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[0\] vssd1 vssd1 vccd1
+ vccd1 _05996_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09169__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__clkinv_4
X_13062_ _07397_ _07400_ _07435_ net889 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a31o_1
XANTENNA__16435__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net280 net2366 net468 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08778__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16821_ net1375 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_8
Xfanout491 _07221_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16752_ net1306 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13964_ net1018 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09341__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ clknet_leaf_118_wb_clk_i _02154_ _00661_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12915_ team_02_WB.instance_to_wrap.top.pc\[14\] _06271_ _02948_ vssd1 vssd1 vccd1
+ vccd1 _02949_ sky130_fd_sc_hd__o21a_1
X_16683_ net1237 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_13895_ net1152 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11932__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ clknet_leaf_26_wb_clk_i _02085_ _00592_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12846_ team_02_WB.instance_to_wrap.top.pc\[28\] _06231_ vssd1 vssd1 vccd1 vccd1
+ _02880_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15565_ clknet_leaf_25_wb_clk_i _02016_ _00523_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _05543_ _05548_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14516_ net1051 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11728_ net340 net2027 net565 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10254__A2 _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ clknet_leaf_56_wb_clk_i _01947_ _00454_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net1129 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11659_ net334 net2031 net572 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09947__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14378_ net1050 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
Xmax_cap603 _05654_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold906 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap614 _04822_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16117_ clknet_leaf_63_wb_clk_i _02563_ _01075_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold917 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold928 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net2326 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _03217_ _03233_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold939 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16048_ clknet_leaf_39_wb_clk_i _02499_ _01006_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08870_ net959 _04303_ _04314_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a32o_1
XANTENNA__09580__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ _03650_ _03653_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15802__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07752_ _03641_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09332__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07683_ _03530_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14719__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15952__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09422_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] net801 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08717__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _05023_ _05027_ _05028_ _05029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[23\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08438__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ _03425_ _04182_ net2719 net938 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__A1 _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09284_ _04955_ _04957_ _04959_ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16640__1211 vssd1 vssd1 vccd1 vccd1 _16640__1211/HI net1211 sky130_fd_sc_hd__conb_1
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08235_ _04089_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1151_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ _04003_ _04026_ _04027_ _04018_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a211o_1
XANTENNA__09938__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07994__C _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15332__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08097_ _03951_ _03956_ _03957_ net225 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__and4_2
XFILLER_0_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout876_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\] net823 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ net401 _06601_ _06413_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11752__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12700_ _06320_ _06325_ _07325_ _04422_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13680_ net1016 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XANTENNA__10484__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10892_ net420 _06536_ _06412_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12631_ _06116_ _06407_ _06455_ net405 net422 vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__a311o_1
X_16816__1370 vssd1 vssd1 vccd1 vccd1 _16816__1370/HI net1370 sky130_fd_sc_hd__conb_1
XFILLER_0_13_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08429__A2 _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10236__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15350_ clknet_leaf_109_wb_clk_i _01801_ _00308_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12562_ net351 net2486 net464 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ net1080 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11513_ _05837_ net432 _07102_ _07111_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[4\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ clknet_leaf_18_wb_clk_i _01732_ _00239_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ net348 net2604 net482 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14232_ net1056 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
X_11444_ _05703_ _05747_ _06013_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__nor3_1
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ net1148 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
X_11375_ net421 _06578_ _06983_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__B1 team_02_WB.instance_to_wrap.top.aluOut\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ _07117_ net228 _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__o21ai_1
X_10326_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\] net851 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__a22o_1
XANTENNA__15825__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ net1114 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ net231 _03060_ _03062_ net890 _03059_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\] net701 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a22o_1
XANTENNA__09905__B _05567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12612__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10188_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\] net832 net756 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\]
+ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16804_ net1358 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
XANTENNA__10132__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14996_ net1172 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
X_13947_ net1045 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
X_16735_ net1289 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08668__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16700__1254 vssd1 vssd1 vccd1 vccd1 _16700__1254/HI net1254 sky130_fd_sc_hd__conb_1
XANTENNA__11662__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15205__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16666_ net1221 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_13878_ net1106 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15617_ clknet_leaf_1_wb_clk_i _02068_ _00575_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12829_ _07377_ _07452_ _07376_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__a21oi_1
X_16597_ clknet_leaf_75_wb_clk_i _02831_ _01470_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13413__A2 _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15548_ clknet_leaf_62_wb_clk_i _01999_ _00506_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09093__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ clknet_leaf_119_wb_clk_i _01930_ _00437_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12493__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08840__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14274__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08020_ _03900_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12924__A1 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold703 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold714 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _05623_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nor2_4
XFILLER_0_110_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11837__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08922_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\] net662 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09553__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net34 net950 _04555_ net2750 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07804_ net341 _03679_ _03672_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08784_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[0\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[0\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__mux2_2
XANTENNA__10042__A _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ _03597_ _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout457_A _06326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1199_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ _03524_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09405_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\] net688 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__a22o_1
XANTENNA__13072__B _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07597_ _03486_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout624_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09336_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] net880 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__a22o_1
XANTENNA__09084__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09267_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] net812 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08831__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07497__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ _04066_ _04097_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15848__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09198_ _04871_ _04873_ _04875_ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ _04003_ _04026_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09792__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _06031_ _06786_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__nor2_1
XANTENNA__11747__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ net462 _05723_ _05769_ net456 net740 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a221o_1
XANTENNA__15998__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11091_ _06248_ net743 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] net443
+ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _05677_ _05700_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__and2_1
Xhold30 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[16\] vssd1 vssd1 vccd1 vccd1
+ net1428 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__B1 _06963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[11\] vssd1 vssd1 vccd1 vccd1
+ net1439 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1161 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
Xhold52 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[0\] vssd1 vssd1 vccd1 vccd1
+ net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[23\] vssd1 vssd1 vccd1 vccd1
+ net1461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15228__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold74 _02601_ vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold85 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[26\] vssd1 vssd1 vccd1
+ vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ net1011 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XANTENNA_input18_A wbm_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12578__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14781_ net1182 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11993_ net1803 net331 net534 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16520_ clknet_leaf_7_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[23\]
+ _01394_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13732_ net1142 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
X_10944_ _06556_ _06557_ _06559_ team_02_WB.instance_to_wrap.top.aluOut\[26\] net460
+ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__o32a_2
XANTENNA__08357__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16451_ clknet_leaf_67_wb_clk_i net1535 _01325_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13663_ net1125 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10875_ _06517_ _06518_ _06520_ team_02_WB.instance_to_wrap.top.aluOut\[28\] net460
+ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__o32a_4
X_15402_ clknet_leaf_51_wb_clk_i _01853_ _00360_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10209__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12614_ _07036_ _07056_ _07076_ _07241_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__and4b_1
X_16382_ clknet_leaf_73_wb_clk_i _02813_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11406__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09075__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net1188 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15333_ clknet_leaf_127_wb_clk_i _01784_ _00291_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12545_ net303 net2242 net466 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08822__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15264_ clknet_leaf_7_wb_clk_i _01715_ _00222_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12476_ net281 net2100 net480 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ net1152 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XANTENNA_5 team_02_WB.instance_to_wrap.top.DUT.read_data2\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11427_ net913 _07032_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__nor2_1
X_15195_ clknet_leaf_119_wb_clk_i _01646_ _00153_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14146_ net1093 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XANTENNA__09783__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _06968_ _06969_ _06970_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[11\]
+ sky130_fd_sc_hd__or3_2
XFILLER_0_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16003__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11657__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\] net736 net688 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a22o_1
X_14077_ net1055 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
X_11289_ team_02_WB.instance_to_wrap.top.pc\[14\] _06334_ vssd1 vssd1 vccd1 vccd1
+ _06907_ sky130_fd_sc_hd__nor2_1
XANTENNA__09535__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ team_02_WB.instance_to_wrap.top.pc\[18\] net943 net942 _03048_ vssd1 vssd1
+ vccd1 vccd1 _01516_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11342__B1 team_02_WB.instance_to_wrap.top.aluOut\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1050 net1053 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__buf_4
Xfanout1061 net1066 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1072 net1077 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1083 net1086 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12488__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14979_ net1041 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07520_ team_02_WB.instance_to_wrap.top.pad.count\[0\] net991 vssd1 vssd1 vccd1 vccd1
+ _03415_ sky130_fd_sc_hd__nand2_1
X_16718_ net1272 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ net1387 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09066__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _04796_ _04798_ _04800_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__or4_4
XFILLER_0_84_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08813__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09052_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\] net786 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10523__A_N _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08003_ _03887_ _03889_ _03892_ _03890_ _03858_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold500 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14732__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold533 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\] net734 net682 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08905_ net978 net910 _04588_ _04589_ _04587_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13067__B net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\] net867 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__a22o_1
Xhold1200 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10136__B2 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout574_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1222 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ net21 net947 net921 net1750 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] vssd1 vssd1 vccd1 vccd1
+ net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1255 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net1583 net957 net926 _04540_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
Xhold1277 team_02_WB.instance_to_wrap.top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 net2675
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12398__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1288 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1299 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07718_ _03581_ _03604_ _03586_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ net745 _04445_ _04449_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__and3_4
XANTENNA__08608__C team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03509_ _03537_ vssd1 vssd1
+ vccd1 vccd1 _03540_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _06227_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09319_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\] net639 _04499_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10591_ team_02_WB.instance_to_wrap.top.pc\[24\] _06241_ vssd1 vssd1 vccd1 vccd1
+ _06243_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08804__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10072__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ net356 net2111 net503 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16026__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net339 net2381 net510 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XANTENNA__13010__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ net1017 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
X_11212_ team_02_WB.instance_to_wrap.top.pc\[15\] _06335_ team_02_WB.instance_to_wrap.top.pc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__a21oi_1
X_12192_ net331 net2505 net518 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11143_ _06184_ _06192_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15050__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15951_ clknet_leaf_33_wb_clk_i _02402_ _00909_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11074_ net437 _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10025_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] net775 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a22o_1
X_14902_ net1186 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
X_15882_ clknet_leaf_44_wb_clk_i _02333_ _00840_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14833_ net1168 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13077__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14764_ net1179 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XANTENNA__12101__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11976_ net2518 net264 net535 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XANTENNA__09296__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08518__C net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ net1148 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
X_16503_ clknet_leaf_129_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[6\]
+ _01377_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10927_ _06363_ _06388_ net390 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__mux2_1
X_14695_ net1166 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11940__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13646_ net1064 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
X_16434_ clknet_leaf_82_wb_clk_i net1521 _01308_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10858_ net385 _06503_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16365_ clknet_leaf_102_wb_clk_i _02798_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13577_ net1170 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
X_10789_ _06434_ _06437_ _06438_ team_02_WB.instance_to_wrap.top.aluOut\[30\] net460
+ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__o32a_4
X_15316_ clknet_leaf_53_wb_clk_i _01767_ _00274_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12528_ net1990 net354 net479 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16296_ clknet_leaf_97_wb_clk_i _02729_ _01239_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15247_ clknet_leaf_31_wb_clk_i _01698_ _00205_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12459_ net337 net2230 net486 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09756__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16519__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ clknet_leaf_46_wb_clk_i _01629_ _00136_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09220__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11387__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14129_ net1029 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout309 _06975_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09508__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15543__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09670_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] net821 net849 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ team_02_WB.instance_to_wrap.top.a1.instruction\[12\] _04407_ _04389_ vssd1
+ vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__o21a_1
X_08552_ net102 net1571 net893 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XANTENNA__12011__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09287__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07503_ net1674 team_02_WB.instance_to_wrap.ramload\[2\] net968 vssd1 vssd1 vccd1
+ vccd1 _02831_ sky130_fd_sc_hd__mux2_1
X_08483_ _04308_ _04309_ net742 net752 net1628 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a32o_1
XANTENNA__11850__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16049__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_A _06834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] net706 net700 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a22o_1
XANTENNA__10054__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] net694 net662 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09747__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold341 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net1750
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A _04468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 _04657_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
Xfanout821 _04638_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_6
Xfanout832 _04678_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09937_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] net819 net766 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\]
+ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__a221o_1
Xfanout843 _04672_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _04655_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
Xfanout865 net868 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_6
Xfanout876 _04668_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_8
Xfanout887 _04374_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
X_09868_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\] net657 net650 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\]
+ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a221o_1
Xhold1030 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_2
Xhold1041 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1052 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ net164 net952 net903 net1549 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1063 team_02_WB.instance_to_wrap.top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 net2461
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\] net783 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1085 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ net355 net2177 net555 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1096 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09278__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11761_ net337 net2204 net561 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XANTENNA__08486__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11760__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03353_ _03354_ vssd1
+ vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__o21a_1
X_10712_ _06359_ _06362_ net365 vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__mux2_1
XANTENNA__10293__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14480_ net1016 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11692_ net332 net2080 net569 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _03310_ _03313_ net1176 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08238__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10643_ _06258_ _06293_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ clknet_leaf_38_wb_clk_i net1539 _01108_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XANTENNA__15416__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input85_A wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ team_02_WB.instance_to_wrap.top.a1.row1\[115\] _03219_ _03223_ team_02_WB.instance_to_wrap.top.a1.row1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a22o_1
X_10574_ team_02_WB.instance_to_wrap.top.pc\[29\] _06225_ vssd1 vssd1 vccd1 vccd1
+ _06226_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15101_ clknet_leaf_116_wb_clk_i _01552_ _00059_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12990__C1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ net295 net2531 net501 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12591__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16081_ clknet_leaf_94_wb_clk_i _02532_ _01039_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[101\]
+ sky130_fd_sc_hd__dfstp_1
X_13293_ _03178_ _03191_ _03182_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__a21o_1
XANTENNA__14372__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ net1166 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09738__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12244_ net272 net2032 net511 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__mux2_1
XANTENNA__09202__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15566__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ net266 net1771 net518 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
X_16653__1220 vssd1 vssd1 vccd1 vccd1 _16653__1220/HI net1220 sky130_fd_sc_hd__conb_1
XANTENNA__10405__A _05175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11126_ _06184_ _06754_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11935__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11057_ net450 _06684_ _06688_ net439 _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a221o_1
X_15934_ clknet_leaf_4_wb_clk_i _02385_ _00892_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07516__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\] net676 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\]
+ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a221o_1
XANTENNA__09910__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15865_ clknet_leaf_107_wb_clk_i _02316_ _00823_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14816_ net1201 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15796_ clknet_leaf_52_wb_clk_i _02247_ _00754_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ net336 net1833 net536 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
XANTENNA__08477__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14747_ net1201 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11670__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14678_ net1196 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16417_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[16\]
+ _01291_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_13629_ net1080 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15096__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10036__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09977__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ clknet_leaf_96_wb_clk_i _02781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11784__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ clknet_leaf_94_wb_clk_i _02712_ _01231_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11536__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07983_ _03834_ _03865_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11845__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _05385_ _05387_ _05388_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09901__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09653_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] net716 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\]
+ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout272_A _06674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__A1 _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ team_02_WB.instance_to_wrap.top.a1.instruction\[5\] _04364_ net910 _04399_
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\] net678 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\]
+ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08535_ net89 net1694 net891 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout537_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1181_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15439__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08466_ _04319_ net1682 _04286_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08483__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08397_ _03411_ _04261_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout704_A _04461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10027__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _04625_ _04698_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10290_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\] net841 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold160 team_02_WB.instance_to_wrap.top.pc\[20\] vssd1 vssd1 vccd1 vccd1 net1558
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _02594_ vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 net128 vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 net137 vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08943__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10750__A1 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _04487_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_8
Xfanout651 _04484_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11755__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 _04480_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
X_13980_ net1123 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
Xfanout673 _04475_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_2
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_4
XANTENNA__09499__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout695 _04467_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_2
X_12931_ _02887_ _02964_ _02888_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15650_ clknet_leaf_46_wb_clk_i _02101_ _00608_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12862_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ net297 net2496 net552 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__mux2_1
X_14601_ net1178 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15581_ clknet_leaf_111_wb_clk_i _02032_ _00539_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12586__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ _05797_ _05836_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10266__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14532_ net1093 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
X_11744_ net271 net2410 net561 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16364__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09671__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ net1132 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
X_11675_ net264 net2586 net570 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__mux2_1
X_16202_ clknet_leaf_37_wb_clk_i _02647_ _01159_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13414_ net2553 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1
+ vccd1 _03299_ sky130_fd_sc_hd__nand2_1
XANTENNA__09959__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _06274_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__or2_1
X_14394_ net1058 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output191_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09423__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ clknet_leaf_6_wb_clk_i net1523 _01091_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13345_ team_02_WB.instance_to_wrap.top.a1.row1\[105\] _03216_ _03239_ team_02_WB.instance_to_wrap.top.a1.row1\[121\]
+ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a22o_1
XANTENNA__11230__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ _04846_ _04866_ _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16064_ clknet_leaf_8_wb_clk_i _02515_ _01022_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13276_ team_02_WB.instance_to_wrap.top.pad.keyCode\[6\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or4b_2
XFILLER_0_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10488_ _04804_ _04823_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__nand2b_1
X_15015_ net1164 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__inv_2
X_12227_ net334 net2346 net512 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10135__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12158_ net328 net2295 net521 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
XANTENNA__11665__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net409 _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__nand2_1
X_12089_ net302 net2487 net526 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15917_ clknet_leaf_24_wb_clk_i _02368_ _00875_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15848_ clknet_leaf_18_wb_clk_i _02299_ _00806_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ clknet_leaf_45_wb_clk_i _02230_ _00737_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10257__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ net1672 net938 net920 _04197_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09662__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08251_ _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15731__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10009__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ _04053_ net224 _04065_ _04052_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__B _05481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13040__A1_N _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput221 net221 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1027_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15111__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ _03854_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] net710 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ _03786_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09636_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net801 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\]
+ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09567_ _05235_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__and2b_1
XANTENNA__13434__B1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout919_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net70 net69 net41 net40 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] net634 _05157_ _05170_
+ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09653__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ net960 _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11460_ _06897_ _07062_ net395 vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09405__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ _06060_ _06063_ net363 vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11391_ net393 _06817_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13130_ team_02_WB.instance_to_wrap.top.a1.nextHex\[1\] team_02_WB.instance_to_wrap.top.a1.nextHex\[2\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[0\] sky130_fd_sc_hd__or2_1
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ _05989_ _05993_ _05994_ _05995_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[0\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13061_ _02946_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__xnor2_1
X_10273_ _05918_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_4
X_12012_ net273 net2178 net468 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
XANTENNA_input48_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16820_ net1374 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15604__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout481 net483 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ net1305 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
Xfanout492 _07220_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963_ net1013 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15702_ clknet_leaf_111_wb_clk_i _02153_ _00660_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12914_ _02909_ _02947_ _02907_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__o21ai_1
X_16682_ net1236 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_13894_ net1139 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09892__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12845_ team_02_WB.instance_to_wrap.top.pc\[28\] _06231_ vssd1 vssd1 vccd1 vccd1
+ _02879_ sky130_fd_sc_hd__and2_1
X_15633_ clknet_leaf_111_wb_clk_i _02084_ _00591_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ clknet_leaf_53_wb_clk_i _02015_ _00522_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12633__D1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _05493_ _05502_ _07398_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ net334 net2406 net564 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ net1127 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XANTENNA__08852__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ clknet_leaf_14_wb_clk_i _01946_ _00453_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14825__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14446_ net1116 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_11658_ net330 net1884 net573 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ team_02_WB.instance_to_wrap.top.pc\[17\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _06261_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14377_ net1025 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
X_11589_ _05999_ _06127_ net446 _07172_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold907 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16116_ clknet_leaf_62_wb_clk_i _02562_ _01074_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12951__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold918 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ net986 net987 _03232_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold929 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15134__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce_dly team_02_WB.instance_to_wrap.top.pad.button_control.debounce
+ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__and2b_2
X_16047_ clknet_leaf_32_wb_clk_i _02498_ _01005_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07820_ _03658_ _03704_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10190__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _03580_ _03622_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07682_ _03554_ _03555_ _03558_ net362 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09421_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\] net817 net789 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09352_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] net796 net756 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\]
+ _05013_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a221o_1
XANTENNA__09096__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09635__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ _04170_ _04171_ _04173_ _04180_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\] net681 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08843__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08234_ _04088_ _04090_ _04064_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ _04018_ _04032_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ _03951_ _03956_ net225 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09020__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11902__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08998_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\] net845 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ _03838_ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15777__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10960_ net388 _06419_ _06461_ _06600_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09874__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\] net736 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ net400 _06535_ _06420_ _06413_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _06408_ _06456_ _06495_ net422 vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__a31oi_1
XANTENNA_input102_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09087__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ net354 net2444 net467 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08834__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ _04604_ _07104_ _07109_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__a211o_1
X_14300_ net1098 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15280_ clknet_leaf_36_wb_clk_i _01731_ _00238_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12492_ net338 net2231 net482 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__mux2_1
XANTENNA__15157__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14231_ net1107 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
X_11443_ _07045_ _07046_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14162_ net1081 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
X_11374_ net449 _06984_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10944__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ net231 _03116_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10325_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] net775 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14093_ net1134 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _07440_ _03061_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09011__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] net732 net664 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16552__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12104__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10187_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] net856 net772 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a22o_1
XANTENNA__10413__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16803_ net1357 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
X_14995_ net1171 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__inv_2
XANTENNA__11943__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ net1288 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
X_13946_ net1045 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XANTENNA__09865__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16665_ team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net106
+ sky130_fd_sc_hd__clkbuf_1
X_13877_ net1120 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15616_ clknet_leaf_12_wb_clk_i _02067_ _00574_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09078__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12828_ _07378_ _07451_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16596_ clknet_leaf_75_wb_clk_i net1649 _01469_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09617__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15547_ clknet_leaf_104_wb_clk_i _01998_ _00505_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11424__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ _05094_ _06249_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15478_ clknet_leaf_108_wb_clk_i _01929_ _00436_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1031 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09250__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold715 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold748 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _05625_ _05627_ _05629_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__or4_2
Xhold759 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] net633 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09002__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ net35 net948 net922 net2226 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10163__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ net341 _03679_ _03660_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__a21boi_1
X_08783_ net1595 net957 net926 _04548_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11853__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ _03581_ _03604_ _03596_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07665_ _03509_ _03537_ _03523_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__a21boi_4
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11154__A team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\] net636 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07596_ _03449_ _03480_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__xor2_1
XANTENNA__09608__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09335_ _05006_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__nor2_2
XANTENNA__16425__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09266_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\] net790 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\]
+ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08217_ _04098_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09197_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] net715 net639 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\]
+ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08148_ _04026_ _04027_ _04003_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09241__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ _03959_ _03965_ _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_4
X_10110_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] net615 _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a22o_1
X_11090_ net912 _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _05677_ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nor2_1
XANTENNA__10154__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[22\] vssd1 vssd1 vccd1 vccd1
+ net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[1\] vssd1 vssd1 vccd1 vccd1
+ net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[24\] vssd1 vssd1 vccd1 vccd1
+ net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[14\] vssd1 vssd1 vccd1 vccd1
+ net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[9\] vssd1 vssd1 vccd1 vccd1
+ net1462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11763__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\] vssd1 vssd1 vccd1 vccd1
+ net1473 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ net1096 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
Xhold86 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\] vssd1 vssd1 vccd1 vccd1
+ net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _02605_ vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11992_ net2169 net326 net534 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
X_14780_ net1181 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09847__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ net1071 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
X_10943_ net441 _06561_ _06569_ net451 _06585_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[26\]
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_39_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16450_ clknet_leaf_75_wb_clk_i net1541 _01324_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10874_ _04416_ _06310_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__nor3_1
X_13662_ net1020 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15401_ clknet_leaf_32_wb_clk_i _01852_ _00359_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ _07126_ _07240_ _07145_ _07108_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16381_ clknet_leaf_73_wb_clk_i _02812_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12594__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ net1200 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XANTENNA__08807__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14375__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12544_ net295 net2388 net464 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15332_ clknet_leaf_19_wb_clk_i _01783_ _00290_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12475_ net273 net2543 net482 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__mux2_1
X_15263_ clknet_leaf_8_wb_clk_i _01714_ _00221_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10408__A _05257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14214_ net1092 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_11426_ _06331_ _07031_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__or2_1
XANTENNA_6 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15194_ clknet_leaf_123_wb_clk_i _01645_ _00152_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_54_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11938__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ net1103 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ net429 _06957_ _06958_ net442 vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\] net636 _05961_ vssd1
+ vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21o_1
X_14076_ net1097 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
X_11288_ net429 _06892_ _06906_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[14\]
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13027_ _06781_ _07336_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\] net821 net853 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10145__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__A1 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1044 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_4
XANTENNA__11342__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1051 net1053 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
Xfanout1062 net1066 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1073 net1077 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_4
XANTENNA__11673__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1084 net1086 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_4
XFILLER_0_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1095 net1138 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09299__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14978_ net1044 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16717_ net1271 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
X_13929_ net1011 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XANTENNA__15322__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16648_ net1386 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16579_ clknet_leaf_82_wb_clk_i net1428 _01452_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09120_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\] net689 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15472__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09471__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ _04730_ _04731_ _04732_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _03851_ _03859_ _03884_ _03849_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09223__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold512 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11848__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold545 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold556 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] net730 net637 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08904_ team_02_WB.instance_to_wrap.top.a1.instruction\[12\] _04407_ _04375_ vssd1
+ vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11149__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__A2 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ net750 _05545_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout1107_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net22 net947 net921 net1730 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1245 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout567_A _07195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[9\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[9\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__mux2_2
Xhold1278 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1289 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
X_07717_ _03606_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or2_1
X_08697_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\] net630 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout734_A _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07648_ _03509_ _03537_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] vssd1 vssd1
+ vccd1 vccd1 _03539_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08608__D team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07579_ _03455_ _03466_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a21bo_2
XANTENNA_fanout901_A _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09318_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] net671 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a22o_1
X_10590_ _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__inv_2
XANTENNA__09462__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] net694 net659 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ net335 net2350 net510 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11211_ net321 net2398 net585 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12191_ net327 net2615 net518 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07537__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _06769_ _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__nand2_1
XANTENNA__13258__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11059__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15950_ clknet_leaf_33_wb_clk_i _02401_ _00908_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11073_ _06704_ _06705_ net409 vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A wbm_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] net857 net797 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\]
+ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a221o_1
X_14901_ net1171 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15881_ clknet_leaf_32_wb_clk_i _02332_ _00839_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12589__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14832_ net1168 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14763_ net1178 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11975_ net1718 net258 net532 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_16502_ clknet_leaf_0_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[5\]
+ _01376_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13714_ net1084 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ net421 _06568_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor2_1
XANTENNA__15495__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14694_ net1196 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
X_16433_ clknet_leaf_82_wb_clk_i net1465 _01307_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13645_ net1130 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
X_10857_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ clknet_leaf_102_wb_clk_i _02797_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net744 net458 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ net444 vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__a221o_1
X_13576_ net1170 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
XANTENNA__09453__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10063__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ clknet_leaf_126_wb_clk_i _01766_ _00273_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ net2708 net345 net477 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16295_ clknet_leaf_100_wb_clk_i _02728_ _01238_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14833__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15246_ clknet_leaf_33_wb_clk_i _01697_ _00204_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09205__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net336 net2417 net484 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11409_ _05658_ _06168_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__xor2_1
X_15177_ clknet_leaf_31_wb_clk_i _01628_ _00135_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12389_ net312 net1820 net494 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14128_ net1021 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
X_14059_ net1026 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XANTENNA__10118__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ team_02_WB.instance_to_wrap.top.a1.instruction\[12\] _04368_ _04377_ net909
+ _04362_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__a311o_1
XANTENNA__08731__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08606__B_N team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15838__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ net103 net1670 net894 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07502_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net2744 net968 vssd1
+ vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ _04305_ _04306_ net742 net751 net1582 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09692__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15988__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09444__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ _04783_ _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and2b_2
XANTENNA__08798__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\] net684 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\]
+ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1057_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold320 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 net148 vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 team_02_WB.instance_to_wrap.top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net1751
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 _04660_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold386 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] vssd1
+ vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _04657_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] net799 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a22o_1
Xfanout822 _04638_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
Xfanout833 _04677_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout844 _04672_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout855 _04655_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_6
XANTENNA__11306__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout866 net868 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
Xfanout877 _04668_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
X_09867_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] net718 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout851_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12710__B _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout899 _04627_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_4
Xhold1031 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1042 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net175 net951 net902 net1514 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08188__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09798_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] net841 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__a22o_1
Xhold1064 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1086 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1097 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ net2702 net955 net927 _04531_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13822__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11760_ net336 net1733 net560 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XANTENNA__08916__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _06360_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11691_ net329 net2097 net569 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10642_ team_02_WB.instance_to_wrap.top.pc\[19\] _06254_ vssd1 vssd1 vccd1 vccd1
+ _06294_ sky130_fd_sc_hd__xnor2_1
X_13430_ _03300_ _03312_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ team_02_WB.instance_to_wrap.top.a1.row1\[19\] _03222_ _03234_ team_02_WB.instance_to_wrap.top.a1.row2\[19\]
+ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] net930 net590 vssd1
+ vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ clknet_leaf_47_wb_clk_i _01551_ _00058_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ net287 net2022 net501 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16080_ clknet_leaf_37_wb_clk_i _02531_ _01038_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13292_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] _03174_ _03200_ _03201_
+ net995 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__o221a_1
XANTENNA_input78_A wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ net1168 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__inv_2
X_12243_ net276 net2739 net509 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11545__A1 _05863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ net260 net2634 net518 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
XANTENNA__10405__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ _05235_ _06031_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09482__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15933_ clknet_leaf_114_wb_clk_i _02384_ _00891_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11056_ _05073_ net430 _06689_ net436 _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10007_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\] net688 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a22o_1
X_15864_ clknet_leaf_121_wb_clk_i _02315_ _00822_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12112__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ net1201 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15795_ clknet_leaf_124_wb_clk_i _02246_ _00753_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11951__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13732__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14746_ net1182 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
X_11958_ net332 net2544 net538 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09674__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10909_ _06548_ _06549_ _06552_ team_02_WB.instance_to_wrap.top.aluOut\[27\] net460
+ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o32a_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16465__D team_02_WB.instance_to_wrap.top.aluOut\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14677_ net1197 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_11889_ net309 net2597 net547 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16416_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[15\]
+ _01290_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_131_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13628_ net1097 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XANTENNA__09426__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16347_ clknet_leaf_101_wb_clk_i _02780_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13559_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03393_ vssd1
+ vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__or4b_1
XANTENNA__14563__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16278_ clknet_leaf_97_wb_clk_i _02711_ _01230_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15229_ clknet_leaf_114_wb_clk_i _01680_ _00187_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10339__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07982_ _03870_ _03871_ _03866_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15660__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] net863 net802 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\]
+ _05382_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11427__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12022__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09652_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\] net724 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08603_ _04365_ _04368_ _04372_ _04379_ _04397_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a221o_1
X_09583_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] net727 net639 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a22o_1
XANTENNA__16016__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ net90 team_02_WB.START_ADDR_VAL_REG\[26\] net891 vssd1 vssd1 vccd1 vccd1
+ _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09665__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11472__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net961 _04317_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ net2017 net935 net918 _04265_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a22o_1
XANTENNA__09417__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12972__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_A _04627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _04625_ _04698_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11527__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 _02779_ vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 team_02_WB.instance_to_wrap.top.a1.data\[5\] vssd1 vssd1 vccd1 vccd1 net1559
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 net142 vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold183 net139 vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_02_WB.instance_to_wrap.top.pad.button_control.noisy vssd1 vssd1 vccd1
+ vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12721__A team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_6
XANTENNA__10750__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout641 _04487_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09919_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] net670 net650 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a22o_1
Xfanout652 net655 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_8
Xfanout663 _04480_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
Xfanout674 _04475_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_8
Xfanout685 net687 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_8
Xfanout696 net699 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_6
X_12930_ _02890_ _02892_ _02962_ _02889_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12861_ team_02_WB.instance_to_wrap.top.pc\[21\] _06253_ vssd1 vssd1 vccd1 vccd1
+ _02895_ sky130_fd_sc_hd__nor2_1
XANTENNA__11771__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600_ net1178 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
X_11812_ net288 net2149 net552 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15580_ clknet_leaf_61_wb_clk_i _02031_ _00538_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16509__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ _07410_ _07413_ _07415_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__o21a_1
XANTENNA__07550__A team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09120__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ net1071 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
X_11743_ net278 net2349 net562 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14462_ net1023 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XANTENNA__09408__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11674_ net259 net2299 net570 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ clknet_leaf_30_wb_clk_i _02646_ _01158_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10018__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ _04182_ _03297_ _03298_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15533__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ team_02_WB.instance_to_wrap.top.pc\[12\] _06276_ vssd1 vssd1 vccd1 vccd1
+ _06277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14393_ net1063 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16132_ clknet_leaf_71_wb_clk_i _02578_ _01090_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13344_ team_02_WB.instance_to_wrap.top.a1.row1\[113\] _03219_ _03245_ _03248_ vssd1
+ vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a211o_1
X_10556_ _06142_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ clknet_leaf_27_wb_clk_i _02514_ _01021_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _03180_ _03183_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__or3_1
XANTENNA__12107__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10416__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ _04603_ _06055_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11518__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15014_ net1165 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
XANTENNA__15683__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ net331 net2527 net514 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__mux2_1
XANTENNA__11946__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ net311 net2353 net521 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11108_ net402 _06505_ _06738_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__a21oi_1
X_12088_ net292 net1972 net524 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08147__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11247__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15916_ clknet_leaf_43_wb_clk_i _02367_ _00874_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11039_ net273 net1796 net584 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15847_ clknet_leaf_13_wb_clk_i _02298_ _00805_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11681__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15778_ clknet_leaf_49_wb_clk_i _02229_ _00736_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07460__A team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09111__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ net1040 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08250_ _04103_ _04104_ _04119_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08870__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08181_ _04030_ net224 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13401__S _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12017__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_3_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput211 net211 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput222 net222 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XANTENNA__09178__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11856__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10193__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07965_ _03804_ _03855_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__xor2_4
XFILLER_0_138_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09704_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\] net737 net697 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\]
+ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07896_ _03744_ _03775_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__xor2_1
XANTENNA__15406__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09635_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\] net814 net853 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__a22o_1
XANTENNA__09350__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout647_A _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09638__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _05216_ _05234_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ net43 net42 net45 net44 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__or4_1
XANTENNA__15556__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout814_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\] net643 _04500_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08448_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\] net917 vssd1 vssd1 vccd1
+ vccd1 _04306_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08379_ _04237_ _04242_ _04244_ _04239_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12945__B1 _07365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10410_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11390_ _06146_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09810__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] net803 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ _05979_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ _02910_ _02912_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10272_ _05920_ _05922_ _05924_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12011_ net276 net2193 net470 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XANTENNA__11766__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16795__1349 vssd1 vssd1 vccd1 vccd1 _16795__1349/HI net1349 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 _07208_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ net1304 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
Xfanout493 _07220_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ net1036 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09877__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15701_ clknet_leaf_114_wb_clk_i _02152_ _00659_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09341__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11684__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12913_ _02910_ _02946_ _02911_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_79_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16681_ net1235 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__12597__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ net1074 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15632_ clknet_leaf_37_wb_clk_i _02083_ _00590_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12844_ team_02_WB.instance_to_wrap.top.pc\[29\] _06228_ vssd1 vssd1 vccd1 vccd1
+ _02878_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09629__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ clknet_leaf_22_wb_clk_i _02014_ _00521_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05493_ _05502_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514_ net1084 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ net330 net2431 net565 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15494_ clknet_leaf_11_wb_clk_i _01945_ _00452_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11440__A2_N _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14445_ net1133 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11657_ net328 net1950 net573 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12626__A _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08823__B net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ net749 _05723_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__o21a_2
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ net1083 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09801__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11588_ _04603_ _06130_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16115_ clknet_leaf_66_wb_clk_i _02561_ _01073_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13327_ _03397_ _03398_ _03231_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__or3_1
Xhold908 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ _05215_ _05234_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o21a_1
XANTENNA__14841__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16046_ clknet_leaf_40_wb_clk_i _02497_ _01004_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13258_ team_02_WB.instance_to_wrap.ramload\[31\] net982 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[31\] sky130_fd_sc_hd__and2_1
XFILLER_0_0_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11676__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ net265 net1953 net515 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap612_A _05071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10175__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ _03146_ _03172_ _03171_ _03148_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15429__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ _03639_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09868__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09332__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ _03554_ net362 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14288__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09420_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] net878 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a22o_1
XANTENNA__12300__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09351_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] net804 net764 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ _05014_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11978__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ _04170_ _04173_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09282_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\] net697 net669 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08233_ _04107_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10650__A1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout228_A _07336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _04046_ _04047_ _04011_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__and3b_1
XFILLER_0_82_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16204__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08095_ _03970_ _03976_ _03979_ _03980_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1137_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16354__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08997_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] net863 net853 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13104__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ _03813_ _03832_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09323__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _03767_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09618_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\] net696 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a221o_1
XANTENNA__12210__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ net388 _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\] net850 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12560_ net342 net2033 net465 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11511_ _05839_ net454 net446 _05838_ _07106_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ net336 net1746 net480 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ net1111 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11442_ _06120_ _07043_ _07044_ net449 vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ net421 _06568_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__a21oi_1
X_14161_ net1029 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input60_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ net381 _05975_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__or2_1
X_13112_ _07410_ _07413_ _07415_ _03117_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o31a_1
XFILLER_0_123_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14092_ net1005 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] net720 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _07391_ _07392_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_123_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10186_ net972 net750 _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15721__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16802_ net1356 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
XFILLER_0_94_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14994_ net1172 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
Xfanout290 _06727_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16733_ net1287 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
X_13945_ net1062 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16664_ net1398 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XANTENNA__12120__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ net1036 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15615_ clknet_leaf_8_wb_clk_i _02066_ _00573_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12827_ _07380_ _07450_ _07379_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__a21o_1
X_16595_ clknet_leaf_75_wb_clk_i _02829_ _01468_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14836__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ clknet_leaf_120_wb_clk_i _01997_ _00504_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12758_ _07381_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15101__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11709_ net265 net2208 net566 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15477_ clknet_leaf_124_wb_clk_i _01928_ _00435_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12689_ _06714_ _06766_ net417 vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ net1127 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14359_ net1107 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold705 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold716 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15251__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold738 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16029_ clknet_leaf_116_wb_clk_i _02480_ _00987_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_08920_ _04598_ _04603_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__or2_1
XANTENNA__10148__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ net36 net947 net921 net2241 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__o22a_1
XANTENNA__09553__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _03676_ _03688_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08782_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[1\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[1\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07733_ _03573_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _03523_ _03538_ _03550_ _03520_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09403_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] net720 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07595_ _03443_ _03485_ _03484_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout345_A _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12073__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _04994_ _04995_ _05008_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__or4_2
XANTENNA__08816__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16794__1348 vssd1 vssd1 vccd1 vccd1 _16794__1348/HI net1348 sky130_fd_sc_hd__conb_1
XANTENNA__10623__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09265_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] net798 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout512_A _07215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08216_ _04066_ _04097_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] net717 net700 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08147_ team_02_WB.instance_to_wrap.top.a1.row2\[34\] net936 net919 _04032_ vssd1
+ vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08078_ _03929_ _03961_ _03932_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a21boi_2
XANTENNA__09792__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout881_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ net899 _05681_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold10 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[22\] vssd1 vssd1 vccd1 vccd1
+ net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[26\] vssd1 vssd1 vccd1 vccd1
+ net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[31\] vssd1 vssd1 vccd1 vccd1
+ net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold43 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[19\] vssd1 vssd1 vccd1 vccd1
+ net1441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[12\] vssd1 vssd1 vccd1 vccd1
+ net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_02_WB.instance_to_wrap.top.pad.button_control.debounce vssd1 vssd1 vccd1
+ vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_02_WB.instance_to_wrap.top.pc\[9\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15894__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 team_02_WB.instance_to_wrap.top.pc\[5\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net1765 net314 net534 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
Xhold98 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[21\] vssd1 vssd1 vccd1
+ vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13730_ net1088 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10942_ _04910_ net430 net428 _06562_ _06584_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15124__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13661_ net1054 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
X_10873_ _06230_ _06309_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15400_ clknet_leaf_110_wb_clk_i _01851_ _00358_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12612_ net426 _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ clknet_leaf_73_wb_clk_i _02811_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13592_ net1200 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15331_ clknet_leaf_45_wb_clk_i _01782_ _00289_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12543_ net289 net1999 net464 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15274__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15262_ clknet_leaf_12_wb_clk_i _01713_ _00220_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12474_ net277 net2666 net481 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10408__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ net1089 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ team_02_WB.instance_to_wrap.top.pc\[8\] _06330_ vssd1 vssd1 vccd1 vccd1 _07031_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15193_ clknet_leaf_106_wb_clk_i _01644_ _00151_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_7 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14144_ net1082 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11356_ net434 _06963_ _06966_ _06965_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09783__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11590__A2 _07179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\] net676 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__a22o_1
X_14075_ net1060 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XANTENNA__12115__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11287_ net440 _06894_ _06900_ net448 _06905_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__o221a_1
XANTENNA__09535__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ net229 _03045_ _03046_ _07445_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] net837 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_4
XANTENNA__08743__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11954__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1044 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_2
XANTENNA__13735__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10169_ _05819_ _05821_ _05823_ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__or4_2
Xfanout1063 net1066 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1074 net1077 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1099 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__buf_4
XANTENNA__16468__D team_02_WB.instance_to_wrap.top.aluOut\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14977_ net1009 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16716_ net1270 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_13928_ net1096 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16647_ net1385 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ net1071 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13470__A _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16578_ clknet_leaf_82_wb_clk_i net1442 _01451_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15617__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15529_ clknet_leaf_24_wb_clk_i _01980_ _00487_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07482__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\] net794 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\]
+ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08001_ _03849_ _03854_ _03887_ _03889_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__or4b_1
XFILLER_0_41_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold502 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold513 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold524 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09774__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12025__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _05591_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11869__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08903_ team_02_WB.instance_to_wrap.top.a1.instruction\[13\] _03396_ _04391_ vssd1
+ vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__o21ai_1
X_09883_ net462 _04504_ net456 _05546_ net741 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a221o_1
XANTENNA__11864__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net23 net949 net923 net1692 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
Xhold1213 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1235 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1246 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ net1601 net955 net926 _04539_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
XANTENNA__15147__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1279 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
X_07716_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _03581_ _03604_ vssd1 vssd1
+ vccd1 vccd1 _03607_ sky130_fd_sc_hd__and3_1
X_08696_ net748 _04442_ _04445_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07647_ _03509_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07578_ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ _03438_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16542__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12708__B _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09317_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] net699 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\] net707 net619 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a22o_1
XANTENNA__10072__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__B _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09179_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\] net823 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13010__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11210_ net461 team_02_WB.instance_to_wrap.top.aluOut\[17\] _06833_ vssd1 vssd1 vccd1
+ vccd1 _06834_ sky130_fd_sc_hd__o21a_2
X_12190_ net313 net2734 net518 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XANTENNA__09765__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11141_ net417 net448 _06766_ _06759_ net437 vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__o32a_1
XFILLER_0_43_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09517__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _06445_ _06452_ net403 vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__mux2_1
Xinput100 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08725__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] net865 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__a22o_1
X_14900_ net1187 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15880_ clknet_leaf_56_wb_clk_i _02331_ _00838_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08649__A team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A wbm_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ net1168 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XANTENNA__13077__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11088__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14762_ net1177 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11974_ net1885 net255 net533 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ clknet_leaf_1_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[4\]
+ _01375_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13713_ net1078 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
X_10925_ net397 _06566_ _06567_ _06425_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14693_ net1157 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16432_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[31\]
+ _01306_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13644_ net1004 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
X_10856_ _06415_ _06502_ net379 vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16363_ clknet_leaf_102_wb_clk_i _02796_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13575_ net1170 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
X_10787_ net912 _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15314_ clknet_leaf_20_wb_clk_i _01765_ _00272_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ net2029 net349 net477 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
X_16294_ clknet_leaf_96_wb_clk_i _02727_ _01237_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15245_ clknet_leaf_23_wb_clk_i _01696_ _00203_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12457_ net331 net2475 net486 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12634__A _06880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ net328 net1873 net584 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XANTENNA__09756__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15176_ clknet_leaf_55_wb_clk_i _01627_ _00134_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08413__C1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ net310 net2579 net495 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ net1129 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ net907 _06277_ _06952_ _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__a32o_1
XANTENNA__09508__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ net1037 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XANTENNA__11684__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net232 _03030_ _03032_ net890 _03029_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a221o_1
X_16793__1347 vssd1 vssd1 vccd1 vccd1 _16793__1347/HI net1347 sky130_fd_sc_hd__conb_1
XFILLER_0_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08550_ net73 net1695 net892 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16565__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ net1594 team_02_WB.instance_to_wrap.ramload\[4\] net968 vssd1 vssd1 vccd1
+ vccd1 _02833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08481_ _04302_ _04303_ net742 net751 net1630 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13404__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ _04763_ _04782_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nand2_1
XANTENNA__10054__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09033_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] net677 net674 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a22o_1
XANTENNA__11859__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold310 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09747__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold321 team_02_WB.instance_to_wrap.top.a1.row2\[16\] vssd1 vssd1 vccd1 vccd1 net1719
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net1730
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold343 team_02_WB.instance_to_wrap.top.a1.row1\[2\] vssd1 vssd1 vccd1 vccd1 net1741
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold365 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold376 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net804 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_8
Xfanout812 _04657_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
X_09935_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\] net807 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a221o_1
Xfanout823 _04638_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_8
Xfanout834 _04677_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_2
XANTENNA_fanout677_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12503__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _04664_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_6
Xfanout856 _04655_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_6
X_09866_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\] net646 _05529_ vssd1
+ vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1010 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 _04667_ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_8
Xhold1021 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _04363_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_4
XANTENNA__09380__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ net178 net954 net905 net1516 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
Xhold1032 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1054 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] net861 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__a22o_1
Xhold1065 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[18\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[18\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__mux2_1
Xhold1087 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1098 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09132__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08679_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\] net679 net675 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
XANTENNA__15932__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__B _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ _05296_ net369 vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__nand2_1
XANTENNA__10293__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ net312 net2151 net569 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _06261_ _06290_ _06292_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10045__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ team_02_WB.instance_to_wrap.top.a1.row1\[59\] _03226_ _03235_ team_02_WB.instance_to_wrap.top.a1.row2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a22o_1
X_10572_ team_02_WB.instance_to_wrap.top.pc\[30\] _06222_ vssd1 vssd1 vccd1 vccd1
+ _06224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09986__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11769__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ net281 net1930 net502 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13291_ _03183_ _03189_ _03192_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15030_ net1195 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
XANTENNA__09199__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ net264 net2250 net511 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XANTENNA__09738__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15312__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16438__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net255 net2282 net517 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ net297 net2572 net582 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15932_ clknet_leaf_63_wb_clk_i _02383_ _00890_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11055_ _05075_ net452 net445 _05074_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__a22o_1
XANTENNA__10702__A _05175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _05660_ _05662_ _05664_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__or4_2
X_15863_ clknet_leaf_119_wb_clk_i _02314_ _00821_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09910__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14814_ net1201 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15794_ clknet_leaf_15_wb_clk_i _02245_ _00752_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09123__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14745_ net1193 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ net329 net1961 net538 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XANTENNA__08477__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08826__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ _04416_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10284__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15005__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14676_ net1197 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ net299 net1918 net546 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16415_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[14\]
+ _01289_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13627_ net1045 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
X_10839_ net363 _06378_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10036__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16346_ clknet_leaf_102_wb_clk_i net1548 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11233__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and4_1
XANTENNA__09977__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11679__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16481__D team_02_WB.instance_to_wrap.top.aluOut\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12509_ net2011 net281 net476 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ clknet_leaf_95_wb_clk_i _02710_ _01229_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13489_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ _03345_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15228_ clknet_leaf_61_wb_clk_i _01679_ _00186_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08937__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11536__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ clknet_leaf_119_wb_clk_i _01610_ _00117_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15805__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ _03827_ _03867_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09720_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] net854 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ _05383_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a221o_1
XANTENNA__12303__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09362__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\] net736 net676 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\]
+ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a221o_1
XANTENNA__12709__A_N _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08602_ _04375_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__nor2_1
XANTENNA__15955__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09582_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] net714 net707 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\]
+ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09114__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ net91 net2671 net894 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10488__A_N _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11472__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\] net917 vssd1 vssd1 vccd1
+ vccd1 _04318_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08395_ _04256_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1167_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10027__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15335__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ net580 _04698_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout794_A _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08928__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[17\] vssd1 vssd1 vccd1
+ vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold151 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[1\] vssd1 vssd1 vccd1
+ vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold162 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[23\] vssd1 vssd1 vccd1
+ vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_02_WB.START_ADDR_VAL_REG\[8\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_02_WB.instance_to_wrap.top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1 net1582
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_02_WB.START_ADDR_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12721__B team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 _04495_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_8
Xfanout631 _04492_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_8
X_09918_ _05574_ _05576_ _05578_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__or4_1
Xfanout642 _04487_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_8
Xfanout653 net655 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12213__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 net667 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_8
Xfanout675 _04475_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_8
X_09849_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] net852 net840 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a22o_1
Xfanout697 net699 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ team_02_WB.instance_to_wrap.top.pc\[21\] _06253_ vssd1 vssd1 vccd1 vccd1
+ _02894_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09105__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ net279 net2290 net552 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12791_ _07409_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08646__B team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14530_ net1090 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
X_11742_ net264 net2648 net563 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XANTENNA__10266__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14461_ net1105 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
X_11673_ net256 net2502 net570 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16200_ clknet_leaf_28_wb_clk_i _02645_ _01157_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13412_ net1486 _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nor2_1
XANTENNA_input90_A wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net750 _04507_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__o21a_2
XFILLER_0_10_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09959__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14392_ net1056 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16792__1346 vssd1 vssd1 vccd1 vccd1 _16792__1346/HI net1346 sky130_fd_sc_hd__conb_1
XFILLER_0_10_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16131_ clknet_leaf_71_wb_clk_i _02577_ _01089_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ team_02_WB.instance_to_wrap.top.a1.row2\[41\] _03230_ _03235_ team_02_WB.instance_to_wrap.top.a1.row2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10555_ _04889_ _04909_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16062_ clknet_leaf_5_wb_clk_i _02513_ _01020_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15828__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ _03184_ _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__nor2_1
X_10486_ _04603_ _06055_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15013_ net1162 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__inv_2
XANTENNA__12715__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ net326 net2294 net514 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09592__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net309 net1828 net523 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15978__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ net394 _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__and2_1
XANTENNA__12123__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net284 net1863 net525 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
XANTENNA__08147__A1 team_02_WB.instance_to_wrap.top.a1.row2\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11038_ net460 team_02_WB.instance_to_wrap.top.aluOut\[23\] _06670_ _06673_ vssd1
+ vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__o22a_2
X_15915_ clknet_leaf_20_wb_clk_i _02366_ _00873_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14839__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15846_ clknet_leaf_12_wb_clk_i _02297_ _00804_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16476__D team_02_WB.instance_to_wrap.top.aluOut\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _06642_ _07335_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__or2_1
X_15777_ clknet_leaf_1_wb_clk_i _02228_ _00735_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10257__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14728_ net1042 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15358__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ net1034 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16603__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10009__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _04043_ _04062_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16329_ clknet_leaf_100_wb_clk_i _02762_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput212 net212 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput223 net223 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09583__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ _03779_ _03805_ _03824_ _03826_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and4b_2
XANTENNA__12033__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\] net684 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a22o_1
X_07895_ _03784_ _03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11872__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] net861 net817 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\]
+ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16133__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07651__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ _05196_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout542_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16739__1293 vssd1 vssd1 vccd1 vccd1 _16739__1293/HI net1293 sky130_fd_sc_hd__conb_1
XANTENNA__11173__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ net104 net71 net105 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__and3_1
XANTENNA__10248__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] net730 net679 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08447_ team_02_WB.instance_to_wrap.top.a1.data\[5\] net915 vssd1 vssd1 vccd1 vccd1
+ _04305_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout807_A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold120_A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08378_ _04249_ _04250_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] net811 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\]
+ _05980_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13828__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\] net724 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\]
+ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a221o_1
XANTENNA__09574__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net266 net1901 net470 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10184__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 _04582_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09326__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 _07226_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ net1011 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 _07223_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout494 _07220_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11782__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ clknet_leaf_46_wb_clk_i _02151_ _00658_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13563__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ team_02_WB.instance_to_wrap.top.pc\[11\] _05548_ _02945_ vssd1 vssd1 vccd1
+ vccd1 _02946_ sky130_fd_sc_hd__a21o_1
X_16680_ net1234 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ net1093 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12843_ team_02_WB.instance_to_wrap.top.pc\[30\] _06225_ vssd1 vssd1 vccd1 vccd1
+ _02877_ sky130_fd_sc_hd__nand2_1
X_15631_ clknet_leaf_32_wb_clk_i _02082_ _00589_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15500__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ clknet_leaf_45_wb_clk_i _02013_ _00520_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10239__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12774_ net750 _04504_ _06220_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14513_ net1079 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ net326 net2703 net565 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
X_15493_ clknet_leaf_127_wb_clk_i _01944_ _00451_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08852__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ net1004 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11656_ net311 net2046 net573 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XANTENNA__15650__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07500__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__B _06688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ net929 _05769_ _06220_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__a21o_1
X_14375_ net1136 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11587_ _05999_ _07172_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__and2_1
XANTENNA__12118__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16114_ clknet_leaf_67_wb_clk_i _02560_ _01072_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap606 _05611_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_2
X_13326_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] net985 _03206_ vssd1 vssd1
+ vccd1 vccd1 _03232_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold909 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ _05238_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16006__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ clknet_leaf_24_wb_clk_i _02496_ _01003_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13257_ net1893 net982 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[30\]
+ sky130_fd_sc_hd__and2_1
X_10469_ net379 _06075_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ net260 net1978 net514 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__mux2_1
X_13188_ _03144_ _02782_ _02781_ _02780_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ net250 net2251 net522 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16156__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11692__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07680_ _03560_ _03566_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07471__A team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15180__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15829_ clknet_leaf_115_wb_clk_i _02280_ _00787_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09350_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] net768 _05024_ _05026_
+ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__a211o_1
XANTENNA__09096__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08301_ _04168_ _04174_ _04176_ _04166_ _04178_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09281_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] net737 _04958_ vssd1
+ vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08843__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ _04113_ _04114_ _04096_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nor3b_1
XANTENNA__09398__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ _04046_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12028__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08094_ _03979_ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11867__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1032_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09556__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09020__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout492_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08996_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] net865 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09308__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _03836_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12698__S _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15523__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16791__1345 vssd1 vssd1 vccd1 vccd1 _16791__1345/HI net1345 sky130_fd_sc_hd__conb_1
XANTENNA_fanout757_A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _03685_ _03727_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_138_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09617_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\] net724 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout924_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] net870 net790 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\]
+ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09087__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _05147_ _05149_ _05151_ _05152_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[20\]
+ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08834__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11510_ net426 _07108_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ net331 net2402 net482 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16029__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09101__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11441_ net412 net438 _06658_ net454 _05703_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10929__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14160_ net1003 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ net406 _06981_ _06982_ net408 vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08940__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13111_ net889 _07416_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__nor2_1
XANTENNA__11777__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14091_ net1024 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13343__A1 team_02_WB.instance_to_wrap.top.a1.row2\[41\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__A team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _02906_ _02950_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ net897 _05889_ _05907_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09011__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10185_ net462 _05795_ _05841_ net456 net740 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16801_ net1355 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
X_14993_ net1172 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
Xfanout280 _06699_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_1
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
X_16732_ net1286 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
XANTENNA__12401__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ net1057 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XANTENNA__10710__A _05296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16663_ net1397 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
X_13875_ net1144 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15614_ clknet_leaf_4_wb_clk_i _02065_ _00572_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12826_ _07382_ _07449_ _07383_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16594_ clknet_leaf_67_wb_clk_i net1430 _01467_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09078__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15545_ clknet_leaf_107_wb_clk_i _01996_ _00503_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12757_ _05094_ _06249_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__nand2_1
XANTENNA__08286__B1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10093__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11708_ net259 net1923 net567 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
X_15476_ clknet_leaf_51_wb_clk_i _01927_ _00434_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ _07026_ _07067_ _07292_ _07141_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__or4b_1
XFILLER_0_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ net1048 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13031__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ net254 net1779 net574 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09786__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14358_ net1109 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XANTENNA__09250__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 team_02_WB.instance_to_wrap.top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1
+ net2115 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11687__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13309_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__or3_1
Xhold728 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14289_ net1078 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
Xhold739 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09538__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07466__A team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16028_ clknet_leaf_48_wb_clk_i _02479_ _00986_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_16738__1292 vssd1 vssd1 vccd1 vccd1 _16738__1292/HI net1292 sky130_fd_sc_hd__conb_1
XANTENNA__09002__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15546__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net37 net949 net923 net2678 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07801_ _03689_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nor2_1
XANTENNA__08761__B2 _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08781_ net1570 net956 net926 _04547_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13407__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _03554_ _03555_ _03568_ _03558_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12311__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15696__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07663_ _03548_ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\] net704 net664 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\]
+ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ _03470_ _03471_ _03451_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] net706 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ _05009_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout240_A _06348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08816__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09264_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] net872 _04942_ vssd1
+ vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _04066_ _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\] net667 _04874_ vssd1
+ vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a21o_1
XANTENNA__13022__B1 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout505_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15076__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09777__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _04003_ _04026_ _04027_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__a21o_2
XANTENNA__11033__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11597__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08077_ _03962_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09529__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16471__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[9\] vssd1 vssd1 vccd1 vccd1
+ net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[6\] vssd1 vssd1 vccd1 vccd1
+ net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[8\] vssd1 vssd1 vccd1 vccd1
+ net1431 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] net882 _04635_ _04644_
+ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__and4_4
Xhold44 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[15\] vssd1 vssd1 vccd1 vccd1
+ net1442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[28\] vssd1 vssd1 vccd1 vccd1
+ net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_02_WB.instance_to_wrap.top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 net1464
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12221__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\] vssd1 vssd1 vccd1 vccd1
+ net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net2312 net309 net535 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
Xhold88 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\] vssd1 vssd1 vccd1 vccd1
+ net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09701__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10941_ net439 _06577_ _06579_ _06580_ _06582_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ net1097 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
X_10872_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net744 net458 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ net444 vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ _06155_ _07178_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ net1198 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08807__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15330_ clknet_leaf_47_wb_clk_i _01781_ _00288_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10075__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ net280 net2048 net465 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09480__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15261_ clknet_leaf_113_wb_clk_i _01712_ _00219_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12473_ net263 net2529 net483 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14212_ net1141 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11424_ _05656_ net432 _07017_ _07030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[8\]
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09768__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15192_ clknet_leaf_122_wb_clk_i _01643_ _00150_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14143_ net1112 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11355_ _05524_ net433 net446 _05522_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] net732 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\]
+ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a221o_1
X_14074_ net1045 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11286_ net434 _06901_ _06902_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__o211a_1
X_13025_ _07387_ _07389_ _07444_ net889 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] net861 net797 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_4
XANTENNA__08743__B2 _04528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_4
XANTENNA__09940__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1053 net1067 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
X_10168_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\] net738 net661 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\]
+ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__a221o_1
Xfanout1064 net1066 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__buf_4
Xfanout1075 net1077 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_4
Xfanout1086 net1138 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
XANTENNA__12131__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__buf_4
XANTENNA__09299__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ _05751_ _05753_ _05755_ _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or4_2
X_14976_ net1009 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_63_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16715_ net1269 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_13927_ net1135 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11970__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16646_ net1384 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13858_ net1091 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16484__D team_02_WB.instance_to_wrap.top.aluOut\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12809_ _07401_ _07402_ _07432_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16577_ clknet_leaf_81_wb_clk_i net1451 _01450_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13789_ net1080 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XANTENNA__10066__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15528_ clknet_leaf_56_wb_clk_i _01979_ _00486_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09471__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13004__B1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15459_ clknet_leaf_43_wb_clk_i _01910_ _00417_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_16669__1224 vssd1 vssd1 vccd1 vccd1 _16669__1224/HI net1224 sky130_fd_sc_hd__conb_1
XFILLER_0_26_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08000_ _03851_ _03856_ _03860_ _03854_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09759__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16790__1344 vssd1 vssd1 vccd1 vccd1 _16790__1344/HI net1344 sky130_fd_sc_hd__conb_1
XFILLER_0_5_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold503 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold514 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12306__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold525 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold536 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold547 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold558 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04627_ _05593_ _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o21ai_1
Xhold569 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11318__B1 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _04379_ _04410_ _04371_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13926__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] _04425_ _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08833_ net24 net947 net921 net1700 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__o22a_1
XANTENNA__07924__A team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1203 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1236 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12041__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10350__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[10\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[10\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_2
Xhold1258 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ _03581_ _03604_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1
+ vccd1 vccd1 _03606_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ net748 _04445_ _04454_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11880__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ _03523_ _03532_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a211o_2
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07577_ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] _03458_ vssd1 vssd1 vccd1
+ vccd1 _03468_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout622_A _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _04991_ _04992_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__and2b_1
XANTENNA__09998__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09462__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\] net682 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__A _05247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09178_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] net870 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09214__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08129_ _03987_ _04010_ _04007_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12216__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ net436 _06765_ _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15861__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11071_ net407 _06455_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput101 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07834__A team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] net845 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12765__A_N _05257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16217__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__B team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1188 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A wbm_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11973_ net1745 net252 net533 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14761_ net1181 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
XANTENNA__11790__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16500_ clknet_leaf_36_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[3\]
+ _01374_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13712_ net1016 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ net580 net379 _06565_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or3b_1
X_14692_ net1163 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15241__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16367__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16431_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[30\]
+ _01305_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__inv_2
X_13643_ net1013 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
X_16737__1291 vssd1 vssd1 vccd1 vccd1 _16737__1291/HI net1291 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ net1186 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16362_ clknet_leaf_102_wb_clk_i _02795_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10786_ _06345_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09453__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12525_ net2495 net338 net477 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
X_15313_ clknet_leaf_19_wb_clk_i _01764_ _00271_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16293_ clknet_leaf_96_wb_clk_i _02726_ _01236_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11260__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15244_ clknet_leaf_53_wb_clk_i _01695_ _00202_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12456_ net328 net2438 net486 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XANTENNA__09205__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ net459 team_02_WB.instance_to_wrap.top.aluOut\[9\] _07014_ _06887_ vssd1
+ vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__o22a_2
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15175_ clknet_leaf_114_wb_clk_i _01626_ _00133_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10435__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12126__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ net300 net2297 net494 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
XANTENNA__10220__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ net1114 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11338_ team_02_WB.instance_to_wrap.top.pc\[12\] _06276_ vssd1 vssd1 vccd1 vccd1
+ _06952_ sky130_fd_sc_hd__or2_1
XANTENNA__11965__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ net1012 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11269_ net914 _06888_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__nor2_1
X_13008_ _07449_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__xor2_1
XANTENNA__09913__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14959_ net1000 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07500_ team_02_WB.instance_to_wrap.top.a1.instruction\[5\] net1781 net968 vssd1
+ vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__mux2_1
XANTENNA__10287__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _04299_ _04300_ net742 net751 net1543 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a32o_1
XANTENNA__09692__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16629_ net1377 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_92_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15734__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09444__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ _04763_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09032_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\] net710 net706 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\]
+ _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15884__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 team_02_WB.instance_to_wrap.top.a1.row1\[0\] vssd1 vssd1 vccd1 vccd1 net1698
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold311 team_02_WB.instance_to_wrap.top.a1.row2\[1\] vssd1 vssd1 vccd1 vccd1 net1709
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 team_02_WB.instance_to_wrap.wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net1720
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold333 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold344 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold366 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 team_02_WB.instance_to_wrap.ramload\[12\] vssd1 vssd1 vccd1 vccd1 net1786
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net804 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
X_09934_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\] net859 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a22o_1
Xhold399 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_8
Xfanout824 _04638_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 _04677_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_8
Xfanout846 _04664_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input8_A wbm_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\] net698 net686 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a22o_1
Xfanout857 _04652_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_8
Xhold1000 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 _04646_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout572_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout879 _04667_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
Xhold1011 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net179 net952 net903 net1509 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
Xhold1033 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15264__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1055 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net1681 net956 net925 _04530_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
Xhold1077 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ net745 _04443_ _04454_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__and3_4
XFILLER_0_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09683__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07629_ _03518_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nor2_2
XFILLER_0_90_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ _06258_ _06291_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08657__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ net271 net2103 net502 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ _03178_ _03182_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ net259 net2234 net509 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10202__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net253 net1974 net517 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10753__A1 _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__A0 _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13566__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net459 team_02_WB.instance_to_wrap.top.aluOut\[20\] _06752_ vssd1 vssd1 vccd1
+ vccd1 _06753_ sky130_fd_sc_hd__o21a_4
XFILLER_0_124_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07564__A team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ clknet_leaf_105_wb_clk_i _02382_ _00889_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11054_ net416 _06682_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10005_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\] net656 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\]
+ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a221o_1
X_15862_ clknet_leaf_112_wb_clk_i _02313_ _00820_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16668__1223 vssd1 vssd1 vccd1 vccd1 _16668__1223/HI net1223 sky130_fd_sc_hd__conb_1
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14813_ net1201 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_15793_ clknet_leaf_17_wb_clk_i _02244_ _00751_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15757__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10269__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14744_ net1194 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11956_ net312 net2637 net538 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09674__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07503__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13207__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ _06308_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__xnor2_1
X_14675_ net1197 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11887_ net292 net2720 net544 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[13\]
+ _01288_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ net1045 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
X_10838_ _06483_ _06484_ net390 vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09426__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16345_ clknet_4_10__leaf_wb_clk_i _02778_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13557_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__or4_1
X_10769_ _04625_ net389 vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__A2 _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ net1946 net272 net478 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__mux2_1
X_13488_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] _03345_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a21o_1
X_16276_ clknet_leaf_94_wb_clk_i _02709_ _01228_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15227_ clknet_leaf_104_wb_clk_i _01678_ _00185_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12439_ net258 net2360 net485 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14860__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13391__C1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ clknet_leaf_109_wb_clk_i _01609_ _00116_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11695__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14109_ net1031 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
X_07980_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03867_ _03868_ vssd1 vssd1
+ vccd1 vccd1 _03870_ sky130_fd_sc_hd__or3_1
X_15089_ clknet_leaf_18_wb_clk_i _01540_ _00047_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15287__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16532__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09650_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\] net672 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08601_ net973 net976 _04385_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\] net699 net671 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08532_ net92 net1632 net892 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09665__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ team_02_WB.instance_to_wrap.top.a1.data\[1\] net915 vssd1 vssd1 vccd1 vccd1
+ _04317_ sky130_fd_sc_hd__or2_1
XANTENNA__11472__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08394_ _03411_ _04261_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1062_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09015_ net580 _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16062__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold130 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[6\] vssd1 vssd1 vccd1
+ vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _02596_ vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09050__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 _02580_ vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 _02602_ vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold174 team_02_WB.instance_to_wrap.top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1 net1572
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 net151 vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16736__1290 vssd1 vssd1 vccd1 vccd1 _16736__1290/HI net1290 sky130_fd_sc_hd__conb_1
Xfanout621 _04495_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12721__C team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09917_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] net718 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a221o_1
Xfanout632 net635 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_8
Xfanout643 _04487_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout954_A _04340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout665 net667 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_4
Xfanout676 net679 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_8
X_09848_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] net812 net791 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\]
+ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a221o_1
Xfanout687 _04470_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_4
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\] net714 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ net271 net1976 net554 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05843_ _05883_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09656__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net258 net2447 net562 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11672_ net252 net1861 net570 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__mux2_1
X_14460_ net1097 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XANTENNA__09408__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ net931 _04504_ _06220_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a21o_1
X_13411_ net1488 _04197_ net828 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
X_14391_ net1107 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16130_ clknet_leaf_66_wb_clk_i _02576_ _01088_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07559__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13342_ team_02_WB.instance_to_wrap.top.a1.row2\[17\] _03234_ _03240_ team_02_WB.instance_to_wrap.top.a1.row2\[9\]
+ _03246_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__a221o_1
XANTENNA_input83_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10554_ _04913_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__or4b_2
X_16061_ clknet_leaf_111_wb_clk_i _02512_ _01019_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10485_ _06120_ _06125_ _06137_ _06119_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a211o_1
X_15012_ net1158 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12224_ net313 net2408 net514 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16555__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12155_ net300 net2318 net520 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__mux2_1
XANTENNA__12404__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _06632_ _06736_ net384 vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__mux2_1
X_12086_ net269 net2243 net524 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
X_15914_ clknet_leaf_46_wb_clk_i _02365_ _00872_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11037_ net909 _06671_ _06672_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and3_1
XANTENNA__11151__A1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A1_N net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15845_ clknet_leaf_126_wb_clk_i _02296_ _00803_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15016__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15776_ clknet_leaf_8_wb_clk_i _02227_ _00734_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ net229 _03014_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14727_ net1042 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11939_ net255 net1971 net537 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09949__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ net1047 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16492__D team_02_WB.instance_to_wrap.top.aluOut\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13609_ net1024 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14589_ net1200 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07469__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16328_ clknet_leaf_80_wb_clk_i _02761_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09280__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16259_ clknet_leaf_94_wb_clk_i _02697_ _01216_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput213 net213 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09032__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12314__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07963_ _03798_ _03852_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] net717 net641 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a221o_1
X_07894_ _03755_ _03757_ _03741_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09886__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net805 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _05216_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _04339_ _04342_ _04344_ net1498 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08846__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _05162_ _05164_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__or4_4
XANTENNA__15302__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08446_ _04304_ net1616 net827 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ _04242_ _04244_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15452__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12945__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09810__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16667__1222 vssd1 vssd1 vccd1 vccd1 _16667__1222/HI net1222 sky130_fd_sc_hd__conb_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09023__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] net728 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16649__1387 vssd1 vssd1 vccd1 vccd1 net1387 _16649__1387/LO sky130_fd_sc_hd__conb_1
XANTENNA__12224__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10252__B team_02_WB.instance_to_wrap.top.DUT.read_data2\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _04605_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 _06131_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ net1100 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _07226_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_4
Xfanout484 _07222_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_8
Xfanout495 _07220_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_4
XANTENNA__09877__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ _02913_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13891_ net1020 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ clknet_leaf_42_wb_clk_i _02081_ _00588_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12842_ team_02_WB.instance_to_wrap.top.pc\[30\] _06225_ vssd1 vssd1 vccd1 vccd1
+ _02876_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09629__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15561_ clknet_leaf_31_wb_clk_i _02012_ _00519_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08837__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12773_ _05461_ _06276_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14512_ net1016 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ net311 net1996 net565 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ clknet_leaf_54_wb_clk_i _01943_ _00450_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11655_ net308 net2133 net575 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
X_14443_ net1013 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12626__C _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ team_02_WB.instance_to_wrap.top.pc\[18\] _06257_ vssd1 vssd1 vccd1 vccd1
+ _06258_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14374_ net1140 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
X_11586_ net423 _06850_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08604__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16113_ clknet_leaf_67_wb_clk_i _02559_ _01071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13325_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net985 vssd1 vssd1 vccd1
+ vccd1 _03231_ sky130_fd_sc_hd__nand2b_1
X_10537_ _06185_ _06189_ _06187_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15945__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16044_ clknet_leaf_53_wb_clk_i _02495_ _01002_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13256_ net2748 net981 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[29\]
+ sky130_fd_sc_hd__and2_1
X_10468_ _04602_ _06055_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12207_ net254 net2073 net513 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux2_1
X_13187_ _03146_ _03170_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__nor2_1
XANTENNA__12134__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10175__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ net246 net1790 net522 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11973__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12069_ _07192_ _07205_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09868__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16487__D team_02_WB.instance_to_wrap.top.aluOut\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15325__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15828_ clknet_leaf_51_wb_clk_i _02279_ _00786_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08828__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15759_ clknet_leaf_33_wb_clk_i _02210_ _00717_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_08300_ _04177_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09280_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\] net700 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15475__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ _04086_ _04108_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12309__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08162_ _04024_ _04032_ _04014_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ _03947_ net225 _03949_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09005__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11449__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10166__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11363__B2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net883 _04648_ _04651_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__and3_4
XANTENNA__11883__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _03820_ net262 _03822_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _03728_ _03729_ _03757_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout652_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1300_A team_02_WB.START_ADDR_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09616_ _05279_ _05281_ _05283_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or4_4
XFILLER_0_35_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] net846 net774 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a22o_1
XANTENNA__08819__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout917_A _04277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] net809 net781 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ _05139_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08429_ net960 _04285_ _04291_ _04292_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12219__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _05702_ _06135_ net432 _05701_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13040__B2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11371_ net395 _06791_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__or2_1
XANTENNA__12743__A _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ net381 _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _02928_ _02931_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14090_ net1014 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13041_ _06888_ net228 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ net897 _05889_ _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_2
X_10184_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] net615 _05840_ vssd1
+ vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a21o_1
XANTENNA__15348__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11793__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16800_ net1354 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
X_16759__1313 vssd1 vssd1 vccd1 vccd1 _16759__1313/HI net1313 sky130_fd_sc_hd__conb_1
X_14992_ net1175 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
Xfanout270 _06891_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_1
Xfanout281 _06699_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
X_16731_ net1285 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
Xfanout292 _06935_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13943_ net1108 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10710__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16662_ net1396 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ net1082 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
X_15613_ clknet_leaf_114_wb_clk_i _02064_ _00571_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12825_ _05135_ _06253_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__a21oi_1
X_16593_ clknet_leaf_65_wb_clk_i net1417 _01466_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15544_ clknet_leaf_122_wb_clk_i _01995_ _00502_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12756_ _05052_ _06246_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07511__S _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ net256 net2172 net566 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15475_ clknet_leaf_125_wb_clk_i _01926_ _00433_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12129__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10438__A _05461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ _07100_ _07314_ _07125_ _07085_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16715__1269 vssd1 vssd1 vccd1 vccd1 _16715__1269/HI net1269 sky130_fd_sc_hd__conb_1
XFILLER_0_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ net1062 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XANTENNA__12909__A2 _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09235__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11638_ net251 net2058 net574 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14357_ net1115 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11569_ _05978_ _06127_ net446 _05977_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold718 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13308_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net985 vssd1 vssd1 vccd1
+ vccd1 _03214_ sky130_fd_sc_hd__nand2_1
Xhold729 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ net1006 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11269__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ clknet_leaf_106_wb_clk_i _02478_ _00985_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13239_ team_02_WB.instance_to_wrap.ramload\[12\] net983 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[12\] sky130_fd_sc_hd__and2_1
XFILLER_0_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10148__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07800_ _03676_ _03688_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nor2_1
X_08780_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[2\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[2\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07731_ _03581_ _03596_ _03600_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07662_ _03551_ _03552_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16666__1221 vssd1 vssd1 vccd1 vccd1 _16666__1221/HI net1221 sky130_fd_sc_hd__conb_1
XFILLER_0_1_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09401_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] net708 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07593_ _03470_ _03471_ _03452_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09332_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net730 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16648__1386 vssd1 vssd1 vccd1 vccd1 net1386 _16648__1386/LO sky130_fd_sc_hd__conb_1
XFILLER_0_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09474__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09263_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] net879 net875 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a22o_1
XANTENNA__12039__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ _04089_ _04090_ _04072_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__a21boi_4
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09194_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] net722 net675 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a22o_1
XANTENNA__09226__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13022__B2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11878__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _04003_ _04026_ _04027_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11033__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1142_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _03917_ _03919_ _03963_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16616__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11336__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11336__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[20\] vssd1 vssd1 vccd1 vccd1
+ net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[27\] vssd1 vssd1 vccd1 vccd1
+ net1421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ _04649_ _04653_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__nor2_1
Xhold34 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[2\] vssd1 vssd1 vccd1 vccd1
+ net1432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08488__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold45 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[10\] vssd1 vssd1 vccd1 vccd1
+ net1443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[15\] vssd1 vssd1 vccd1 vccd1
+ net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_02_WB.instance_to_wrap.top.pc\[0\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _03817_ _03818_ _03813_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a21o_1
XANTENNA__12836__A1 _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\] vssd1 vssd1 vccd1 vccd1
+ net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold89 team_02_WB.instance_to_wrap.top.pc\[31\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ net420 _06133_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10871_ net911 _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15790__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ _06054_ _06349_ _06561_ _07237_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input100_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ net1168 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XANTENNA__09465__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12541_ net272 net2460 net466 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ clknet_leaf_63_wb_clk_i _01711_ _00218_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16146__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ net260 net2194 net483 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__mux2_1
XANTENNA__09217__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14211_ net1020 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XANTENNA__11788__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11423_ net442 _07019_ _07026_ net449 _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15191_ clknet_leaf_118_wb_clk_i _01642_ _00149_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11575__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07567__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14142_ net1022 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11354_ net415 _06056_ _06531_ _06147_ net455 vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] net716 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a22o_1
X_14073_ net1061 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11285_ _05399_ net433 _06903_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13024_ _02955_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__xnor2_1
X_10236_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] net773 net761 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output152_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 net1015 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 net1023 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_4
XANTENNA__08743__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12412__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\] net726 net637 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a22o_1
Xfanout1032 net1067 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_2
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1054 net1057 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_4
Xfanout1065 net1066 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
XFILLER_0_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_2
Xfanout1087 net1095 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_4
X_14975_ net1007 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
X_10098_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] net718 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a221o_1
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_2
X_16714_ net1268 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
X_13926_ net1139 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16645_ net1216 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ net1146 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12808_ _07404_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__or2_1
XANTENNA__09456__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16576_ clknet_leaf_81_wb_clk_i net1401 _01449_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13788_ net1123 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15527_ clknet_leaf_14_wb_clk_i _01978_ _00485_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12739_ team_02_WB.instance_to_wrap.top.i_ready net988 vssd1 vssd1 vccd1 vccd1 _07363_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14863__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15458_ clknet_leaf_49_wb_clk_i _01909_ _00416_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13004__B2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11698__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ net1025 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ clknet_leaf_112_wb_clk_i _01840_ _00347_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold504 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold526 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold559 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net899 net605 vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08901_ _04365_ _04368_ _04379_ _04397_ _04360_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a311o_1
X_09881_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] net615 _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08832_ net25 net949 net923 net2278 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
XANTENNA__12322__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1204 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 net110 vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ net1598 net957 net925 _04538_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
Xhold1248 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16019__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10350__B _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1259 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ _03581_ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08694_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\] net647 net643 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a221o_1
XANTENNA__09695__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07645_ _03497_ _03528_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A _06132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ _03455_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ _04972_ _04990_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] net728 net726 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16758__1312 vssd1 vssd1 vccd1 vccd1 _16758__1312/HI net1312 sky130_fd_sc_hd__conb_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11006__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09586__B _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\] net790 net754 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _03971_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__xor2_2
XFILLER_0_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10525__B _05481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08059_ _03945_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__nand2_1
X_11070_ _06144_ _06196_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12740__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_10021_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] net805 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a22o_1
XANTENNA__12232__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__A _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16714__1268 vssd1 vssd1 vccd1 vccd1 _16714__1268/HI net1268 sky130_fd_sc_hd__conb_1
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14760_ net1177 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
X_11972_ net2042 net248 net533 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08946__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ net1129 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
X_10923_ net388 _06416_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11493__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14691_ net1196 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ clknet_leaf_68_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[29\]
+ _01304_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13642_ net1054 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10854_ _06367_ _06371_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16361_ clknet_leaf_101_wb_clk_i _02794_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13573_ net1170 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__inv_2
X_10785_ team_02_WB.instance_to_wrap.top.pc\[29\] _06344_ team_02_WB.instance_to_wrap.top.pc\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15312_ clknet_leaf_37_wb_clk_i _01763_ _00270_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12524_ net1865 net336 net476 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16292_ clknet_leaf_97_wb_clk_i _02725_ _01235_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ clknet_leaf_20_wb_clk_i _01694_ _00201_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12455_ net314 net2550 net486 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12407__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__A _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ team_02_WB.instance_to_wrap.top.pc\[9\] net907 _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\]
+ _07013_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__a221o_1
X_15174_ clknet_leaf_3_wb_clk_i _01625_ _00132_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ net291 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net492 vssd1
+ vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ net1131 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11337_ net426 _06937_ _06951_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[12\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_123_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14056_ net1098 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
X_11268_ team_02_WB.instance_to_wrap.top.pc\[15\] _06335_ vssd1 vssd1 vccd1 vccd1
+ _06888_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16647__1385 vssd1 vssd1 vccd1 vccd1 net1385 _16647__1385/LO sky130_fd_sc_hd__conb_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _07381_ _07383_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nand2_1
X_10219_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\] net647 net627 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a22o_1
XANTENNA__12142__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11199_ _06028_ net431 net447 _05276_ _06583_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09017__A _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14858__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11981__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ net1001 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09677__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16495__D team_02_WB.instance_to_wrap.top.aluOut\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13909_ net1119 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14889_ net1187 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16628_ net1376 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09429__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16559_ clknet_leaf_29_wb_clk_i net1453 _01432_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_09100_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[29\] net593 vssd1
+ vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09031_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] net729 net697 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12317__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09601__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 team_02_WB.instance_to_wrap.top.a1.row2\[10\] vssd1 vssd1 vccd1 vccd1 net1699
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold312 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold323 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold334 team_02_WB.instance_to_wrap.top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1 net1732
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold345 team_02_WB.instance_to_wrap.top.a1.row1\[3\] vssd1 vssd1 vccd1 vccd1 net1743
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold378 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] net867 net775 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a22o_1
Xhold389 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_6
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08530__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout814 net816 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout825 _04557_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A _05863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 _04677_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_4
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] net673 net637 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\]
+ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__a221o_1
XANTENNA__12052__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout847 _04664_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_8
Xfanout858 _04652_ vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15409__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 _04642_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_8
Xhold1012 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net180 net951 net902 net1477 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
XANTENNA__09380__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 team_02_WB.instance_to_wrap.top.pad.keyCode\[5\] vssd1 vssd1 vccd1 vccd1
+ net2432 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _05451_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__nor2_4
Xhold1045 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11891__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_A _07195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1056 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[19\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[19\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__mux2_1
Xhold1078 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09132__A2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08677_ net745 _04442_ _04445_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__and3_1
XANTENNA__12672__C1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ _03483_ _03506_ _03487_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03444_ _03445_ vssd1 vssd1
+ vccd1 vccd1 _03450_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12975__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net931 net590 vssd1
+ vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_106_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09840__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ _04908_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[26\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__12227__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12240_ net254 net1819 net510 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
XANTENNA__09199__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ net246 net1927 net517 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12751__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11122_ net908 _06751_ _06750_ _06749_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold890 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
X_15930_ clknet_leaf_121_wb_clk_i _02381_ _00888_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11053_ net422 _06687_ _06686_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a21oi_2
XANTENNA__15089__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] net728 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ clknet_leaf_116_wb_clk_i _02312_ _00819_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14812_ net1201 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XANTENNA__13582__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ clknet_leaf_39_wb_clk_i _02243_ _00750_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09659__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09123__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ net1194 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
X_11955_ net309 net2285 net539 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _06232_ _06233_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__and2b_1
X_14674_ net1196 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11886_ net285 net2356 net544 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16413_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[12\]
+ _01287_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ net1062 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _06362_ _06384_ net365 vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16344_ clknet_leaf_100_wb_clk_i _02777_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13556_ net1532 _03391_ net884 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__o21a_1
XANTENNA__09831__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ net580 net379 vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__or2_1
X_12507_ net1712 net276 net478 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12137__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16275_ clknet_leaf_94_wb_clk_i _02708_ _01227_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_13487_ net2061 _03345_ _03346_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a21oi_1
X_10699_ _05094_ net372 vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__nand2_1
X_15226_ clknet_leaf_116_wb_clk_i _01677_ _00184_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12438_ net256 net2154 net486 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08937__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15157_ clknet_leaf_115_wb_clk_i _01608_ _00115_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12369_ net243 net1944 net492 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14108_ net1085 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15088_ clknet_leaf_28_wb_clk_i _01539_ _00046_ vssd1 vssd1 vccd1 vccd1 team_02_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ net1111 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10181__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09362__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16757__1311 vssd1 vssd1 vccd1 vccd1 _16757__1311/HI net1311 sky130_fd_sc_hd__conb_1
XFILLER_0_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08600_ _04380_ _04389_ _04391_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and3_1
XANTENNA__15701__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\] net711 net647 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\]
+ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a221o_1
XANTENNA__09114__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08531_ net93 net1567 net892 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08462_ _04316_ net1741 net827 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08393_ net2008 net935 net918 _04263_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09822__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16207__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16713__1267 vssd1 vssd1 vccd1 vccd1 _16713__1267/HI net1267 sky130_fd_sc_hd__conb_1
XANTENNA__10356__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[31\] net592 vssd1
+ vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_66_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13382__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1 net1518
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13667__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold131 _02585_ vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10196__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold142 team_02_WB.instance_to_wrap.top.a1.data\[0\] vssd1 vssd1 vccd1 vccd1 net1540
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 team_02_WB.instance_to_wrap.top.a1.data\[1\] vssd1 vssd1 vccd1 vccd1 net1551
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold164 team_02_WB.instance_to_wrap.top.a1.data\[2\] vssd1 vssd1 vccd1 vccd1 net1562
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 net127 vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 net149 vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout682_A _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 net131 vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09916_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] net705 net693 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout622 _04495_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
Xfanout633 net635 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09889__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout644 _04486_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_6
Xfanout655 _04483_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09880__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_8
X_09847_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] net864 net860 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a22o_1
Xfanout677 net679 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_4
Xfanout688 _04468_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15381__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 _04463_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12510__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09778_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] net650 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ _05443_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09105__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ net1610 net955 net924 _04521_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A1 _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11740_ net255 net2134 net562 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10120__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ net249 net2620 net570 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__mux2_1
XANTENNA__12746__A _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16646__1384 vssd1 vssd1 vccd1 vccd1 net1384 _16646__1384/LO sky130_fd_sc_hd__conb_1
XFILLER_0_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ net1492 _04215_ net828 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10622_ _06272_ _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nand2_1
X_14390_ net1109 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09813__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10423__A1 _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13341_ team_02_WB.instance_to_wrap.top.a1.row1\[57\] _03226_ _03237_ team_02_WB.instance_to_wrap.top.a1.row2\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ _04932_ _04951_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__o21bai_1
X_16060_ clknet_leaf_63_wb_clk_i _02511_ _01018_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13272_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[5\] team_02_WB.instance_to_wrap.top.pad.keyCode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__or4b_2
XANTENNA_input76_A wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10484_ _04699_ net430 _06133_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15011_ net1151 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11796__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ net309 net2471 net515 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__mux2_1
XANTENNA__13577__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10187__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09592__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net294 net2293 net520 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15724__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11105_ _06678_ _06735_ net377 vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12085_ net325 net2119 net524 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09344__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15913_ clknet_leaf_24_wb_clk_i _02364_ _00871_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11036_ _06244_ _06245_ _06302_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15844_ clknet_leaf_55_wb_clk_i _02295_ _00802_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13428__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15775_ clknet_leaf_10_wb_clk_i _02226_ _00733_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _02964_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ net1042 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11938_ net250 net2088 net537 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12778__A_N _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14657_ net1043 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
X_11869_ net239 net2660 net545 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ net1089 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588_ net1181 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16327_ clknet_leaf_92_wb_clk_i _02760_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13539_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\]
+ _03377_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14871__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16258_ clknet_leaf_94_wb_clk_i _02696_ _01215_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
X_15209_ clknet_leaf_24_wb_clk_i _01660_ _00167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_16189_ clknet_leaf_66_wb_clk_i _02635_ _01147_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
Xoutput214 net214 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10904__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09583__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13116__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07962_ _03798_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\] net645 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a22o_1
X_07893_ _03741_ _03755_ _03757_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09632_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] net781 net761 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ _05299_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a221o_1
XANTENNA__12330__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09563_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[18\] net592 vssd1
+ vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08514_ team_02_WB.instance_to_wrap.wb.curr_state\[0\] net957 _04343_ vssd1 vssd1
+ vccd1 vccd1 _04344_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09494_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\] net718 net675 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ _05160_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__a221o_1
XANTENNA__10102__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10653__A1 team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08445_ net960 _04302_ _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout430_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1172_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout528_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08376_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04228_ vssd1 vssd1 vccd1
+ vccd1 _04249_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15747__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12505__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09574__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11381__A2 _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 net433 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09326__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 _04436_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _07226_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 _07222_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ team_02_WB.instance_to_wrap.top.pc\[10\] _05593_ _02943_ vssd1 vssd1 vccd1
+ vccd1 _02944_ sky130_fd_sc_hd__a21o_1
Xfanout496 net499 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_6
XANTENNA__12240__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13890_ net1088 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10341__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08657__C team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12841_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10892__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13860__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15560_ clknet_leaf_86_wb_clk_i _02011_ _00518_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12772_ _05421_ _06271_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ net1127 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
X_11723_ net308 net2663 net567 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XANTENNA__10644__A1 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15491_ clknet_leaf_43_wb_clk_i _01942_ _00449_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15277__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1037 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
X_11654_ net299 net1840 net573 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XANTENNA__16522__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10605_ net749 _05679_ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__o21a_2
XFILLER_0_68_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08065__A2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14373_ net1087 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
X_11585_ net398 _07022_ _07175_ net411 vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ clknet_leaf_66_wb_clk_i _02558_ _01070_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_16756__1310 vssd1 vssd1 vccd1 vccd1 _16756__1310/HI net1310 sky130_fd_sc_hd__conb_1
X_13324_ net986 net987 _03208_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10536_ _05297_ _05315_ _05318_ _06183_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap608 _05480_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16043_ clknet_leaf_21_wb_clk_i _02494_ _01001_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ net1666 net981 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[28\]
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09014__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12415__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _04602_ _06055_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07509__S _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ net253 net1748 net513 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13186_ _02782_ _03162_ _02783_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _04785_ _06050_ _04783_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12137_ net244 net2399 net522 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09317__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ net233 net1894 net530 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12150__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ _06038_ net430 net445 _05032_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16712__1266 vssd1 vssd1 vccd1 vccd1 _16712__1266/HI net1266 sky130_fd_sc_hd__conb_1
XANTENNA__10332__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15827_ clknet_leaf_124_wb_clk_i _02278_ _00785_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16052__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12085__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15758_ clknet_leaf_40_wb_clk_i _02209_ _00716_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14709_ net1035 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15689_ clknet_leaf_31_wb_clk_i _02140_ _00647_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _04084_ _04109_ _04112_ _04088_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ _04014_ _04024_ _04032_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08092_ _03947_ _03949_ net225 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12325__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09556__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11363__A2 team_02_WB.instance_to_wrap.top.aluOut\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08994_ net882 _04648_ _04651_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__and3_2
XANTENNA__09308__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _03820_ _03822_ net262 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__A2 _06734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12060__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03764_ _03765_ _03766_ vssd1
+ vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\] net708 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout645_A _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] net823 net866 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout812_A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] net869 net817 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\]
+ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10809__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ team_02_WB.instance_to_wrap.top.a1.row1\[18\] net827 vssd1 vssd1 vccd1 vccd1
+ _04292_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__A2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _04204_ _04223_ _04232_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11051__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11370_ _06896_ _06980_ net386 vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ _05965_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nor2_8
XFILLER_0_63_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ _07366_ _03058_ team_02_WB.instance_to_wrap.top.pc\[16\] net944 vssd1 vssd1
+ vccd1 vccd1 _01514_ sky130_fd_sc_hd__a2bb2o_1
X_10252_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[2\] vssd1 vssd1 vccd1
+ vccd1 _05907_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08014__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10183_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] _04367_ _04426_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a22o_1
Xfanout1203 net1204 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08949__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ net1175 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__inv_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
Xfanout271 _06674_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout282 _06699_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_1
X_16730_ net1284 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
X_13942_ net1108 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
Xfanout293 _06935_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10314__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09180__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ net1395 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13873_ net1028 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ clknet_leaf_61_wb_clk_i _02063_ _00570_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13590__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _07386_ _07447_ _07384_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__a21oi_1
X_16592_ clknet_leaf_66_wb_clk_i net1402 _01465_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ clknet_leaf_118_wb_clk_i _01994_ _00501_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12755_ _05053_ _06246_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10719__A _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15912__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07494__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11706_ net250 net2413 net566 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15474_ clknet_leaf_26_wb_clk_i _01925_ _00432_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _06946_ _06964_ _07006_ _07044_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10438__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14425_ net1064 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11637_ net248 net2288 net574 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14356_ net1038 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XANTENNA__09786__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ _06112_ _06155_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ net985 net987 _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__nor3b_1
Xhold708 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__inv_2
Xhold719 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ net1127 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XANTENNA__12145__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ net403 _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16026_ clknet_leaf_116_wb_clk_i _02477_ _00984_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13238_ net1713 net982 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[11\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09538__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11984__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _03150_ _03154_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16498__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _03614_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09171__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire613_A _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16568__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07661_ _03516_ _03545_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09400_ _05073_ _05074_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and2b_2
XFILLER_0_1_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07592_ _03477_ _03478_ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\] net719 _05000_ _05007_
+ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _04934_ _04936_ _04938_ _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08213_ _04048_ _04095_ _04094_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09193_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\] net711 net694 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\]
+ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout226_A _07336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11033__A1 _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _04016_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nand2_1
XANTENNA__09777__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ _03920_ _03923_ _03953_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__or3_1
XANTENNA__12055__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1135_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09529__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[11\] vssd1 vssd1 vccd1 vccd1
+ net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[28\] vssd1 vssd1 vccd1 vccd1
+ net1422 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _04656_ net886 _04637_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__and3b_4
XANTENNA_fanout762_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[23\] vssd1 vssd1 vccd1 vccd1
+ net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[16\] vssd1 vssd1 vccd1 vccd1
+ net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07928_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__inv_2
Xhold57 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[12\] vssd1 vssd1 vccd1 vccd1
+ net1455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_02_WB.instance_to_wrap.top.pc\[14\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold79 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[5\] vssd1 vssd1 vccd1
+ vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09701__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15935__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ _06344_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] net674 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07476__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12540_ net275 net2694 net466 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__mux2_1
XANTENNA__10075__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12471_ net256 net2598 net481 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
XANTENNA__12754__A _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ net1090 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ _06120_ _07025_ _07027_ net438 _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15190_ clknet_leaf_109_wb_clk_i _01641_ _00148_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16711__1265 vssd1 vssd1 vccd1 vccd1 _16711__1265/HI net1265 sky130_fd_sc_hd__conb_1
XANTENNA__10232__C1 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ net1054 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
X_11353_ net414 _06540_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10274__A _05928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net728 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14072_ net1055 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11284_ _05402_ net455 net446 _05401_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__a22o_1
XANTENNA__13585__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ _02900_ _02901_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__nor2_1
X_10235_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\] net865 net781 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\]
+ _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10535__B1 _05193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15465__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 net1015 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1011 net1015 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1022 net1023 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_4
XANTENNA__08304__A1_N _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_4
XANTENNA__09940__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\] net698 _05822_ vssd1
+ vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a21o_1
Xfanout1044 net1049 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1055 net1057 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
XFILLER_0_83_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1077 net1138 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_2
Xfanout1088 net1095 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
X_14974_ net1007 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
X_10097_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] net730 net698 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09153__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1099 net1104 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16713_ net1267 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
X_13925_ net1074 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16644_ net1215 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
X_13856_ net1075 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12807_ _05633_ _05636_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ net1045 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XANTENNA__10449__A _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16575_ clknet_leaf_81_wb_clk_i net1452 _01448_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10999_ _04991_ net430 _06630_ _06636_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__a221o_1
XANTENNA__10066__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12738_ team_02_WB.instance_to_wrap.top.a1.state\[0\] _07359_ _07361_ _07362_ vssd1
+ vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__o22a_1
X_15526_ clknet_leaf_12_wb_clk_i _01977_ _00484_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15457_ clknet_leaf_2_wb_clk_i _01908_ _00415_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12669_ _07005_ _07065_ _07130_ _07146_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__and4_1
XFILLER_0_115_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14408_ net1096 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XANTENNA__09759__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15388_ clknet_leaf_63_wb_clk_i _01839_ _00346_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14339_ net1068 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold505 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold516 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold527 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold538 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
X_16659__1393 vssd1 vssd1 vccd1 vccd1 net1393 _16659__1393/LO sky130_fd_sc_hd__conb_1
XANTENNA__11318__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16009_ clknet_leaf_24_wb_clk_i _02460_ _00967_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_08900_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09880_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08831_ net26 net947 net921 net1683 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o22a_1
XANTENNA__09931__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1205 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1216 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[11\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[11\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__mux2_2
Xhold1238 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1249 team_02_WB.instance_to_wrap.top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 net2647
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ _03596_ _03600_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08693_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\] net639 net635 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07644_ _03508_ _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03460_ _03461_ _03463_ vssd1
+ vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout343_A _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _04972_ _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__nor2_1
XANTENNA__10057__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09998__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11889__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15338__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] net739 net722 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\]
+ _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout510_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09176_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\] net831 _04856_ vssd1
+ vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08127_ _03978_ _03981_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08058_ _03903_ _03942_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__xor2_2
XFILLER_0_43_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12513__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10020_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net749 _05680_ vssd1
+ vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__o21a_2
XANTENNA__09383__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput103 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09922__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11971_ net2467 net242 net533 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12749__A _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ net1062 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XANTENNA__08946__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ net385 _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__nand2_1
XANTENNA__11493__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10296__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14690_ net1166 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16113__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13641_ net1011 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
X_10853_ net408 _06495_ _06498_ _06499_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10048__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16360_ clknet_leaf_101_wb_clk_i _02793_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12442__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ net1186 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__inv_2
X_10784_ _06224_ _06226_ _06313_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__o31a_1
XFILLER_0_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15311_ clknet_leaf_33_wb_clk_i _01762_ _00269_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11799__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12523_ net2252 net330 net477 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__mux2_1
X_16291_ clknet_leaf_96_wb_clk_i _02724_ _01234_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15242_ clknet_leaf_51_wb_clk_i _01693_ _00200_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12454_ net309 net2201 net487 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10716__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11405_ net913 _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15173_ clknet_leaf_127_wb_clk_i _01624_ _00131_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12385_ net286 net1917 net493 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14124_ net1005 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10220__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11336_ net440 _06939_ _06945_ net435 _06950_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14055_ net1156 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11267_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] net826 _06321_ _04583_ vssd1
+ vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__a31o_4
XANTENNA__10732__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09374__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ _02896_ _02960_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__xnor2_1
X_10218_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] net715 net667 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a221o_1
XANTENNA__09913__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11198_ net417 _06822_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11039__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] net807 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a221o_1
XANTENNA__09017__B _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09126__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14957_ net1002 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13908_ net1052 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10287__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14888_ net1186 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16627_ net1206 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13839_ net1124 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XANTENNA__16606__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16558_ clknet_leaf_36_wb_clk_i net1421 _01431_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ clknet_leaf_115_wb_clk_i _01960_ _00467_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ clknet_leaf_64_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[24\] _01363_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] net713 net633 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\]
+ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15630__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11539__A2 team_02_WB.instance_to_wrap.top.aluOut\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 team_02_WB.instance_to_wrap.ramload\[25\] vssd1 vssd1 vccd1 vccd1 net1700
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold324 team_02_WB.START_ADDR_VAL_REG\[30\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_02_WB.instance_to_wrap.top.a1.row2\[8\] vssd1 vssd1 vccd1 vccd1 net1755
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15780__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\] net763 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a221o_1
Xhold368 team_02_WB.instance_to_wrap.top.a1.row1\[56\] vssd1 vssd1 vccd1 vccd1 net1766
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold379 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12333__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10642__A team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 _04659_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_6
XANTENNA__09365__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] net702 net692 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout837 _04676_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_8
Xfanout848 _04664_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_A _06935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _04652_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08814_ net181 net951 net902 net1528 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
Xhold1002 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1
+ net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _05453_ _05455_ _05457_ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__or4_1
Xhold1035 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09117__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net1599 net955 net924 _04529_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a22o_1
Xhold1057 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout460_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1079 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710__1264 vssd1 vssd1 vccd1 vccd1 _16710__1264/HI net1264 sky130_fd_sc_hd__conb_1
XFILLER_0_75_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08676_ _04452_ _04460_ _04465_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ _03483_ _03487_ _03506_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__and3_2
XANTENNA__12719__D _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_A _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10089__A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07558_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] _03438_ _03442_ _03448_ vssd1
+ vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07489_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] team_02_WB.instance_to_wrap.ramload\[16\]
+ net965 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
XANTENNA__12508__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09228_ _04898_ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__nor2_4
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09159_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\] net710 net665 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10202__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ net245 net2617 net517 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11121_ _06296_ _06297_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12243__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold880 team_02_WB.instance_to_wrap.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net2278
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11052_ net405 _06407_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__or2_1
XANTENNA__13863__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\] net644 _05663_ vssd1
+ vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a21o_1
X_15860_ clknet_leaf_46_wb_clk_i _02311_ _00818_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09108__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A wbm_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ net1203 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
X_15791_ clknet_leaf_31_wb_clk_i _02242_ _00749_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10269__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14742_ net1194 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
X_11954_ net300 net1711 net538 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10905_ _06231_ net744 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] net443
+ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a221o_1
X_14673_ net1193 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13207__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net268 net1998 net544 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16658__1392 vssd1 vssd1 vccd1 vccd1 net1392 _16658__1392/LO sky130_fd_sc_hd__conb_1
XFILLER_0_50_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16412_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[11\]
+ _01286_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13624_ net1054 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10836_ _06355_ _06359_ net364 vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13555_ _03391_ net884 _03390_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__and3b_1
X_16343_ clknet_leaf_100_wb_clk_i _02776_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ net401 _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__nor2_1
XANTENNA__12418__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12506_ net2197 net265 net479 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16274_ clknet_leaf_97_wb_clk_i _02707_ _01226_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13486_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] _03345_ net873 vssd1 vssd1
+ vccd1 vccd1 _03346_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ _04744_ _06051_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16009__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15225_ clknet_leaf_106_wb_clk_i _01676_ _00183_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12437_ net252 net1909 net485 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09595__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15156_ clknet_leaf_53_wb_clk_i _01607_ _00114_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ net237 net2501 net492 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ net1058 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ net459 team_02_WB.instance_to_wrap.top.aluOut\[13\] _06934_ vssd1 vssd1 vccd1
+ vccd1 _06935_ sky130_fd_sc_hd__o21a_4
XFILLER_0_61_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15087_ clknet_leaf_82_wb_clk_i _01538_ _00045_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12153__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net358 net1898 net504 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
XANTENNA__09347__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ net1110 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XANTENNA__10181__B _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13773__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15183__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15989_ clknet_leaf_124_wb_clk_i _02440_ _00947_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_08530_ net95 net1722 net891 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ net960 _04314_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08392_ _04257_ _04258_ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12957__A1 _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07833__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09013_ _04692_ _04695_ _04696_ _04697_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[31\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout306_A _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13382__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 team_02_WB.instance_to_wrap.top.pc\[25\] vssd1 vssd1 vccd1 vccd1 net1508
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[12\] vssd1 vssd1 vccd1
+ vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09050__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[16\] vssd1 vssd1 vccd1
+ vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold143 team_02_WB.instance_to_wrap.top.pc\[17\] vssd1 vssd1 vccd1 vccd1 net1541
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold154 team_02_WB.instance_to_wrap.top.a1.data\[4\] vssd1 vssd1 vccd1 vccd1 net1552
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_02_WB.START_ADDR_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold176 team_02_WB.instance_to_wrap.top.pc\[10\] vssd1 vssd1 vccd1 vccd1 net1574
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 net124 vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13134__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold198 team_02_WB.instance_to_wrap.top.a1.hexop\[1\] vssd1 vssd1 vccd1 vccd1 net1596
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] net642 _05577_ vssd1
+ vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a21o_1
Xfanout623 _04495_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_8
Xfanout645 _04486_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_4
XANTENNA_fanout675_A _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout656 net659 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_8
X_09846_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\] net815 net772 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\]
+ _05505_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a221o_1
Xfanout667 _04478_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_6
Xfanout689 _04468_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09777_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] net726 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout842_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[28\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[28\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15676__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ net747 _04454_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ net244 net2451 net570 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ team_02_WB.instance_to_wrap.top.pc\[13\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _06273_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14019__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13340_ net987 _03244_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10423__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10552_ _06143_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ _03181_ _03182_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__nor2_1
XANTENNA__13858__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10483_ _04703_ net455 net447 _04700_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a22o_1
XANTENNA__12762__A _05175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_129_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15010_ net1151 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09577__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ net301 net1738 net514 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__mux2_1
XANTENNA__16301__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input69_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09041__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12153_ net286 net2556 net522 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _06350_ _06354_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__nand2_1
X_12084_ net319 net1854 net527 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16451__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11035_ _06244_ _06245_ _06302_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__or3_1
X_15912_ clknet_leaf_18_wb_clk_i _02363_ _00870_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12701__S team_02_WB.instance_to_wrap.top.aluOut\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15843_ clknet_leaf_43_wb_clk_i _02294_ _00801_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12986_ _02887_ _02888_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__nand2b_1
X_15774_ clknet_leaf_6_wb_clk_i _02225_ _00732_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__B2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ net1042 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11937_ net246 net2164 net537 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
XANTENNA__08855__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11868_ _04577_ _07188_ _07199_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or3_1
X_14656_ net999 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13607_ net1135 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
X_10819_ net420 _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__nor2_1
XANTENNA__12148__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14587_ net1047 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11799_ net359 net2704 net558 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16326_ clknet_leaf_92_wb_clk_i _02759_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09280__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11987__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13469_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] _03335_ _03336_ vssd1
+ vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16257_ clknet_leaf_92_wb_clk_i _02695_ _01214_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09568__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ clknet_leaf_57_wb_clk_i _01659_ _00166_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
X_16188_ clknet_leaf_66_wb_clk_i _02634_ _01146_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09032__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput215 net215 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15549__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ clknet_leaf_41_wb_clk_i _01590_ _00097_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07961_ _03825_ _03826_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ _05361_ _05363_ _05365_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or4_2
XFILLER_0_78_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07892_ _03772_ _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__and2_1
XANTENNA__15699__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] net845 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09740__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09562_ _05227_ _05231_ _05232_ _05233_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[18\]
+ sky130_fd_sc_hd__or4_4
X_08513_ net988 team_02_WB.instance_to_wrap.wb.curr_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _04343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] net739 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08846__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08444_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\] net917 vssd1 vssd1 vccd1
+ vccd1 _04303_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12058__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand2_1
XANTENNA__13052__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1165_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__S net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1273_A team_02_WB.START_ADDR_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09559__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16657__1391 vssd1 vssd1 vccd1 vccd1 net1391 _16657__1391/LO sky130_fd_sc_hd__conb_1
XFILLER_0_121_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16805__1359 vssd1 vssd1 vccd1 vccd1 _16805__1359/HI net1359 sky130_fd_sc_hd__conb_1
Xfanout420 net424 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout431 net433 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 _04604_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12521__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 _06129_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout464 _07225_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 _07226_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 _07222_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] net715 net623 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a22o_1
Xfanout497 net499 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _04624_ _06316_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12771_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08837__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12757__A _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__B team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14510_ net1117 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
X_11722_ net299 net2121 net565 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
X_15490_ clknet_leaf_50_wb_clk_i _01941_ _00448_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08446__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ net294 net2261 net572 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
X_14441_ net1024 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ net929 _05723_ _06220_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a21o_1
XANTENNA__09798__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14372_ net1146 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
X_11584_ net392 _07096_ _07174_ net404 vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16111_ clknet_leaf_70_wb_clk_i _02557_ _01069_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13323_ _03137_ _03220_ _03228_ _03210_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__or4b_1
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ _05168_ _05174_ _05193_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07586__A team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13254_ net2741 net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[27\]
+ sky130_fd_sc_hd__and2_1
X_16042_ clknet_leaf_44_wb_clk_i _02493_ _01000_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ _06057_ _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__nor2_1
XANTENNA__09014__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ net248 net2626 net513 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12642__D _07269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13185_ _02782_ _03164_ _03169_ _03149_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10397_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08773__B2 _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ net239 net1731 net522 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12067_ net358 net2489 net528 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XANTENNA__12431__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14212__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11018_ _06654_ net413 net436 vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15991__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15826_ clknet_leaf_11_wb_clk_i _02277_ _00784_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15757_ clknet_leaf_43_wb_clk_i _02208_ _00715_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08828__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ team_02_WB.instance_to_wrap.top.pc\[27\] net943 net942 _02998_ vssd1 vssd1
+ vccd1 vccd1 _01525_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ net1042 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XANTENNA__15221__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ clknet_leaf_18_wb_clk_i _02139_ _00646_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14639_ net1194 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14882__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08160_ _04022_ _03978_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09789__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16309_ clknet_leaf_78_wb_clk_i _02742_ _01252_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08091_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__inv_2
XANTENNA__16497__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13337__A1 team_02_WB.instance_to_wrap.top.a1.row2\[40\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13004__A1_N _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08993_ net883 _04644_ _04651_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and3_1
XANTENNA__12341__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _03831_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07875_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03726_ _03756_ vssd1 vssd1
+ vccd1 vccd1 _03766_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\] net644 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09545_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] net854 net778 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout540_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] net861 net878 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ team_02_WB.instance_to_wrap.top.a1.data\[10\] net915 _04290_ vssd1 vssd1
+ vccd1 vccd1 _04291_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13025__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15714__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14792__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _04205_ _04224_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12516__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ _04159_ _04167_ _04144_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ _05967_ _05969_ _05971_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__or4_4
XFILLER_0_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15864__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11339__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _05891_ _05901_ _05904_ _05906_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[2\]
+ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10011__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__B2 _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _05837_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10562__A1 _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_2
XANTENNA__12251__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout250 _06521_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14990_ net1173 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
Xfanout261 _06586_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08507__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _06674_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_1
X_13941_ net1120 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
Xfanout294 _06935_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_1
XANTENNA__11511__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16660_ net1394 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__15244__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ net1016 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15611_ clknet_leaf_105_wb_clk_i _02062_ _00569_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12823_ _07385_ _07446_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__nand2_1
X_16591_ clknet_leaf_65_wb_clk_i net1422 _01464_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10078__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ clknet_leaf_111_wb_clk_i _01993_ _00500_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ _04629_ _05006_ _05011_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10719__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ net246 net2605 net566 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _06569_ _06653_ _07309_ _07312_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__or4_1
XANTENNA__13016__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15473_ clknet_leaf_19_wb_clk_i _01924_ _00431_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ net243 net2157 net574 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
X_14424_ net1054 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XANTENNA__09796__A _05461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09235__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12426__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11567_ _05977_ _06000_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__a21o_1
X_14355_ net1128 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10735__A _05461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10250__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13111__A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13306_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] net986 _03211_ vssd1 vssd1
+ vccd1 vccd1 _03212_ sky130_fd_sc_hd__and3b_1
X_10518_ _05503_ _05521_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__and2b_1
X_14286_ net1116 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11498_ _07021_ _07096_ net386 vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08787__A_N net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ team_02_WB.instance_to_wrap.ramload\[10\] net981 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[10\] sky130_fd_sc_hd__and2_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16025_ clknet_leaf_117_wb_clk_i _02476_ _00983_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10449_ _05677_ net367 vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10002__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09943__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ _02782_ _03153_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10553__A1 _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12119_ net268 net1934 net586 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XANTENNA__12161__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ team_02_WB.instance_to_wrap.top.pc\[6\] net945 net941 _03107_ vssd1 vssd1
+ vccd1 vccd1 _01504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14877__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07660_ _03521_ _03549_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ clknet_leaf_130_wb_clk_i _02260_ _00767_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07591_ _03447_ _03472_ _03480_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a22o_2
XFILLER_0_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ net1343 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_0_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10069__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09330_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] net735 net623 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ _05001_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09474__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\] net859 net804 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\]
+ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16656__1390 vssd1 vssd1 vccd1 vccd1 net1390 _16656__1390/LO sky130_fd_sc_hd__conb_1
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13005__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08682__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16804__1358 vssd1 vssd1 vccd1 vccd1 _16804__1358/HI net1358 sky130_fd_sc_hd__conb_1
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08212_ _04048_ _04077_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09192_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\] net689 net687 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15887__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09226__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11569__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03967_ vssd1 vssd1 vccd1
+ vccd1 _04029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12336__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10241__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08074_ _03930_ _03960_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__xor2_2
XFILLER_0_86_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15117__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13956__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09934__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout588_A _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[17\] vssd1 vssd1 vccd1 vccd1
+ net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15267__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ net883 _04636_ _04648_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold25 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[5\] vssd1 vssd1 vccd1 vccd1
+ net1423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[24\] vssd1 vssd1 vccd1 vccd1
+ net1434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[18\] vssd1 vssd1 vccd1 vccd1
+ net1445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16512__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ _03764_ _03814_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__xor2_1
Xhold58 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[30\] vssd1 vssd1 vccd1 vccd1
+ net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_02_WB.instance_to_wrap.top.pc\[11\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout755_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14787__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07858_ _03706_ _03736_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07789_ net341 _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11415__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09528_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] net717 net713 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\]
+ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ _05126_ _05128_ _05130_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__or4_4
XFILLER_0_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ net250 net2484 net481 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09217__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ _05657_ _06135_ net455 _05658_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11024__A2 _06658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12246__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14140_ net1098 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11352_ net450 _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] net684 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a22o_1
X_14071_ net1112 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ net424 net437 _06408_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _07366_ _03043_ team_02_WB.instance_to_wrap.top.pc\[19\] net944 vssd1 vssd1
+ vccd1 vccd1 _01517_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_input51_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net845 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a22o_1
XANTENNA__09925__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10535__A1 _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1012 net1015 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10165_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] net666 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a22o_1
Xfanout1023 net1032 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_4
Xfanout1045 net1046 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_4
XFILLER_0_41_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_4
Xfanout1067 net5 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
X_14973_ net999 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
X_10096_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\] net646 _05754_ vssd1
+ vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a21o_1
Xfanout1078 net1086 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
Xfanout1089 net1095 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_4
XFILLER_0_136_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16712_ net1266 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13924_ net1143 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16643_ net1214 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_138_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13855_ net1118 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ _07405_ _07428_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o21ai_1
X_16574_ clknet_leaf_91_wb_clk_i net1411 _01447_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13786_ net1038 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XANTENNA__09456__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ _04993_ net452 net445 _04992_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10449__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15525_ clknet_leaf_127_wb_clk_i _01976_ _00483_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12737_ _03423_ _07357_ net961 _03418_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15456_ clknet_leaf_7_wb_clk_i _01907_ _00414_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ _07099_ _07101_ _07084_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14407_ net1152 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12156__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ net294 net2494 net576 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15387_ clknet_leaf_104_wb_clk_i _01838_ _00345_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12599_ net72 net989 _07227_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__mux2_1
XANTENNA__10223__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14338_ net1091 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
Xhold506 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11995__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13776__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold539 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14269_ net1054 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XANTENNA__09916__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16008_ clknet_leaf_56_wb_clk_i _02459_ _00966_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16535__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08589__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08830_ net27 net947 net921 net1666 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__o22a_1
Xhold1206 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net1629 net956 net925 _04537_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1217 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
X_07712_ _03574_ _03576_ _03578_ _03602_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08692_ net748 _04442_ _04443_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and3_1
XANTENNA__14400__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09695__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07643_ _03503_ _03507_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11235__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ _03461_ _03463_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__nand2_1
XANTENNA__09447__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _04626_ team_02_WB.instance_to_wrap.top.DUT.read_data2\[24\] net593 vssd1
+ vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08655__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_A _07055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12855__A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09244_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\] net630 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1078_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08544__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16065__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\] net880 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__a22o_1
XANTENNA__11006__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12066__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__A _05257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_A _07218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10214__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _03993_ _03996_ _03998_ _04000_ _03974_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__o311a_1
XFILLER_0_82_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08057_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03942_ _03943_ vssd1 vssd1
+ vccd1 vccd1 _03945_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout872_A _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__A1 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__B2 _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput104 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XANTENNA__15902__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08959_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ _04632_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_98_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11970_ net2573 net238 net533 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ _06501_ _06563_ net379 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__mux2_1
XANTENNA__11493__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10852_ net403 _06485_ net418 vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__a21oi_1
X_13640_ net1090 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10783_ _04416_ _06314_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__nor2_1
XANTENNA__11245__A2 _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ net1186 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15310_ clknet_leaf_40_wb_clk_i _01761_ _00268_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12522_ net1966 net328 net477 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__mux2_1
X_16290_ clknet_leaf_96_wb_clk_i _02723_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.lcd_rs
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input99_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ clknet_leaf_29_wb_clk_i _01692_ _00199_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ net300 net1899 net486 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11404_ team_02_WB.instance_to_wrap.top.pc\[9\] _06331_ vssd1 vssd1 vccd1 vccd1 _07012_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15432__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15172_ clknet_leaf_55_wb_clk_i _01623_ _00130_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12384_ net267 net2612 net492 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09610__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11335_ net449 _06946_ _06949_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__a21oi_1
X_14123_ net1027 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11266_ _04422_ _06321_ _06324_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21o_2
X_14054_ net1139 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10732__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15582__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\] net691 net643 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a22o_1
X_13005_ _06721_ net226 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ net400 _06601_ _06818_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803__1357 vssd1 vssd1 vccd1 vccd1 _16803__1357/HI net1357 sky130_fd_sc_hd__conb_1
X_10148_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\] net857 net793 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14956_ net1041 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_10079_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] net851 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\]
+ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09677__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09314__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ net1144 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
X_14887_ net1168 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16626_ clknet_leaf_68_wb_clk_i _02860_ _01499_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_13838_ net1116 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XANTENNA__09429__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16557_ clknet_leaf_35_wb_clk_i net1419 _01430_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13769_ net1028 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ clknet_leaf_50_wb_clk_i _01959_ _00466_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12984__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ clknet_leaf_64_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[23\] _01362_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15439_ clknet_leaf_34_wb_clk_i _01890_ _00397_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09062__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09601__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 team_02_WB.instance_to_wrap.top.pc\[30\] vssd1 vssd1 vccd1 vccd1 net1701
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold314 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold325 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15925__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold358 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] net851 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13261__A_N net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout805 _04658_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout816 _04654_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
X_09862_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\] net634 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a221o_1
Xfanout827 _04286_ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
Xfanout838 _04676_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_4
Xfanout849 _04662_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_8
Xhold1003 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ net182 net951 net902 net1501 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
Xhold1014 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\] net670 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\]
+ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1036 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[20\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[20\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1069 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] net686 net682 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ _04469_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15305__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1195_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07626_ _03513_ _03516_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07557_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1 vccd1 _03448_
+ sky130_fd_sc_hd__or3_1
XANTENNA_fanout620_A _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12975__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07488_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] net2379 net964 vssd1
+ vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09227_ _04900_ _04902_ _04904_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] net695 net689 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09053__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ _03994_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09089_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] net850 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a22o_1
XANTENNA__12524__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08800__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _06253_ net743 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] net443
+ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold870 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold881 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ net398 _06396_ _06685_ net411 vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__o211a_1
Xhold892 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08022__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\] net720 net696 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10979__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ net1203 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
X_15790_ clknet_leaf_40_wb_clk_i _02241_ _00748_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09659__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input14_A wbm_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1201 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XANTENNA__11466__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ net293 net2130 net536 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10904_ net911 _06547_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__nor2_1
X_14672_ net1167 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ net324 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\] net544 vssd1
+ vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16411_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[10\]
+ _01285_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ net1111 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
X_10835_ _04826_ _06210_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11603__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16342_ clknet_leaf_100_wb_clk_i _02775_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13554_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\]
+ _03387_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__and3_1
XANTENNA__09292__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ net388 _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09831__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ net1815 net260 net479 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16273_ clknet_leaf_92_wb_clk_i _02706_ _01225_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ net238 net2497 net582 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
X_13485_ _03345_ net873 _03344_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__and3b_1
XFILLER_0_125_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15224_ clknet_leaf_123_wb_clk_i _01675_ _00182_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13376__C1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ net246 net2522 net485 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
XANTENNA__09044__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ clknet_leaf_126_wb_clk_i _01606_ _00113_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12434__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ _04576_ _04578_ _07199_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__or3_4
XFILLER_0_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14106_ net1059 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
X_11318_ _06271_ net743 _06887_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__a211o_1
X_15086_ clknet_leaf_77_wb_clk_i _01537_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_12298_ net351 net2653 net504 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14037_ net1117 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
X_11249_ _06151_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09898__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12103__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15988_ clknet_leaf_46_wb_clk_i _02439_ _00946_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08858__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14939_ net1033 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08460_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\] net917 vssd1 vssd1 vccd1
+ vccd1 _04315_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08883__A team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ clknet_leaf_59_wb_clk_i _02843_ _01482_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08391_ _04257_ _04260_ _04258_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09283__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09822__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] net869 net805 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\]
+ _04682_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09035__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__A0 _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 team_02_WB.instance_to_wrap.busy_o vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13382__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[4\] vssd1 vssd1 vccd1
+ vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12344__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 _02591_ vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10196__A2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 _02595_ vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_02_WB.instance_to_wrap.top.pc\[26\] vssd1 vssd1 vccd1 vccd1 net1542
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold155 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[24\] vssd1 vssd1 vccd1
+ vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold166 team_02_WB.instance_to_wrap.top.a1.data\[11\] vssd1 vssd1 vccd1 vccd1 net1564
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_02_WB.instance_to_wrap.top.a1.data\[8\] vssd1 vssd1 vccd1 vccd1 net1575
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold188 team_02_WB.instance_to_wrap.top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1 net1586
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] net714 net709 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a22o_1
Xhold199 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net1597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1110_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout624 net627 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09889__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 _04489_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout646 _04486_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_6
XANTENNA_input6_A wbm_ack_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\] net836 net760 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__a221o_1
Xfanout657 net659 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_4
XANTENNA_fanout570_A _07193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout668 _04477_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_6
Xfanout679 _04474_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
XANTENNA_fanout668_A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09776_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ net1688 net955 net924 _04520_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08849__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout835_A _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14795__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] _04439_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__and3b_2
XFILLER_0_7_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10120__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07609_ _03467_ _03473_ _03468_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08589_ team_02_WB.instance_to_wrap.top.a1.instruction\[5\] net910 _04385_ vssd1
+ vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12519__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10620_ team_02_WB.instance_to_wrap.top.pc\[13\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _06272_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13070__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13070__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09813__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ _06202_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__or2_1
X_16802__1356 vssd1 vssd1 vccd1 vccd1 _16802__1356/HI net1356 sky130_fd_sc_hd__conb_1
XFILLER_0_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__or4b_2
XANTENNA__08732__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09026__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10482_ _04585_ _04596_ _04603_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__or3_4
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12221_ net291 net2701 net512 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__mux2_1
XANTENNA__12254__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10187__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12152_ net269 net1703 net520 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11103_ net422 _06733_ _06732_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a21oi_2
X_12083_ net318 net2344 net525 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11034_ net911 _06668_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__o21bai_1
X_15911_ clknet_leaf_17_wb_clk_i _02362_ _00869_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15842_ clknet_leaf_50_wb_clk_i _02293_ _00800_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ clknet_leaf_114_wb_clk_i _02224_ _00731_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ net989 net911 _04437_ _06642_ net943 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a41o_1
XFILLER_0_8_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ net1040 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ net243 net2124 net537 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14655_ net1007 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12429__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10738__A _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11867_ net235 net1842 net549 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XANTENNA__15770__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13606_ net1091 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10818_ net396 _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
XANTENNA__09265__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14586_ net1045 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11798_ net351 net2684 net556 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ clknet_leaf_90_wb_clk_i _02758_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_13537_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] _03377_
+ net884 vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10749_ _05836_ net369 vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13349__C1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16256_ clknet_leaf_97_wb_clk_i _02694_ _01213_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] _03335_ net1176 vssd1
+ vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15207_ clknet_leaf_14_wb_clk_i _01658_ _00165_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12419_ net294 net1851 net488 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16187_ clknet_leaf_71_wb_clk_i _02633_ _01145_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12164__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
X_13399_ _03143_ _03271_ _03296_ net1183 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_51_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput216 net216 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
X_15138_ clknet_leaf_51_wb_clk_i _01589_ _00096_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09039__A _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15150__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08791__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _03841_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__nand2_2
X_15069_ clknet_leaf_84_wb_clk_i _01520_ _00032_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07891_ _03780_ _03779_ _03778_ _03750_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_65_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09630_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\] net857 net797 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09561_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\] net879 net875 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ _05218_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08512_ net6 _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09492_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\] net647 net627 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10102__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09502__A _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08443_ team_02_WB.instance_to_wrap.top.a1.data\[6\] net915 vssd1 vssd1 vccd1 vccd1
+ _04302_ sky130_fd_sc_hd__or2_1
XANTENNA__12339__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08374_ _04242_ _04244_ _04240_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09256__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13959__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09008__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12074__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__A2_N _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15643__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 net424 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _06322_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 _07225_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout476 _07224_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ _05486_ _05488_ _05490_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__or4_4
Xfanout487 _07222_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_8
XFILLER_0_96_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10341__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] net853 net845 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12770_ _06271_ _05421_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11721_ net293 net1924 net564 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XANTENNA__12249__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11153__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14440_ net1089 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XANTENNA__09247__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11652_ net283 net2520 net574 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10277__B _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13869__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ net928 _05679_ net590 vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a21o_1
X_14371_ net1069 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ net366 _07136_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12773__A _05461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16110_ clknet_leaf_66_wb_clk_i _02556_ _01068_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input81_A wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13322_ team_02_WB.instance_to_wrap.top.a1.row1\[56\] _03226_ _03227_ team_02_WB.instance_to_wrap.top.a1.row1\[0\]
+ _03224_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ _05257_ _05275_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08462__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ clknet_leaf_24_wb_clk_i _02492_ _00999_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13253_ net2278 net981 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[26\]
+ sky130_fd_sc_hd__and2_1
X_10465_ _06086_ _06117_ net418 vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11357__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ net242 net2561 net512 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ _03150_ _03153_ _03158_ _03148_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__o31a_1
X_10396_ _04824_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12135_ _04576_ _04579_ _07188_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__or3_4
XFILLER_0_23_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12066_ net352 net2248 net528 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ net396 _06123_ _06651_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10332__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15825_ clknet_leaf_18_wb_clk_i _02276_ _00783_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15756_ clknet_leaf_43_wb_clk_i _02207_ _00714_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ net229 _02994_ _02997_ _04362_ _02995_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09486__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14707_ net1035 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11919_ net285 net2114 net542 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XANTENNA__12159__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A _04602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15687_ clknet_leaf_16_wb_clk_i _02138_ _00645_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ team_02_WB.instance_to_wrap.top.pc\[3\] _05889_ _02932_ vssd1 vssd1 vccd1
+ vccd1 _02933_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14638_ net1193 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09238__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13034__B2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14569_ net1011 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11596__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16308_ clknet_leaf_80_wb_clk_i _02741_ _01251_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ _03970_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16239_ clknet_leaf_70_wb_clk_i _00009_ _01196_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09410__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10020__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08992_ net882 _04644_ _04651_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__and3_4
XANTENNA__14403__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07943_ _03832_ _03833_ _03819_ net262 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07874_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03756_ _03726_ vssd1 vssd1
+ vccd1 vccd1 _03765_ sky130_fd_sc_hd__o21ai_1
X_16801__1355 vssd1 vssd1 vccd1 vccd1 _16801__1355/HI net1355 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09613_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] net685 _05282_ vssd1
+ vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a21o_1
XANTENNA__12858__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_A _05956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__A_N _07183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09544_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08547__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11284__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] net777 _05138_ _05148_
+ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout533_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08426_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\] net917 vssd1 vssd1 vccd1
+ vccd1 _04290_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15196__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08357_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04221_ _04228_ vssd1 vssd1
+ vccd1 vccd1 _04232_ sky130_fd_sc_hd__or3b_2
XFILLER_0_50_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ _04162_ _04164_ _04157_ _04161_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12536__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11339__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10250_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] net878 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09401__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10181_ net412 _05836_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1205 net5 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_4
XANTENNA__10562__A2 _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__A1 _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 _06348_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout251 _06521_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_1
Xfanout262 _03826_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_2
X_13940_ net1035 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
Xfanout273 _06674_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10314__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 _06912_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_1
XANTENNA__07715__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout295 _06753_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09180__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13871_ net1125 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15610_ clknet_leaf_120_wb_clk_i _02061_ _00568_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12822_ _05216_ _06257_ _07445_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__a21o_1
X_16590_ clknet_leaf_64_wb_clk_i net1424 _01463_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09468__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15541_ clknet_leaf_114_wb_clk_i _01992_ _00499_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15539__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ _05006_ _05011_ _04629_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14983__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11704_ net244 net2078 net566 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
X_15472_ clknet_leaf_34_wb_clk_i _01923_ _00430_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12684_ _06509_ _06635_ _07310_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ net1114 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ net238 net2584 net574 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11611__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ net1079 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
X_11566_ _05999_ _06155_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__nor2_1
XANTENNA__09640__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10735__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__nor2_1
X_10517_ _05378_ _05398_ _06151_ _05356_ _05337_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__o32a_1
X_14285_ net1131 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11497_ _07060_ _07095_ net380 vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16024_ clknet_leaf_123_wb_clk_i _02475_ _00982_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13236_ team_02_WB.instance_to_wrap.ramload\[9\] net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[9\]
+ sky130_fd_sc_hd__and2_1
X_10448_ _06093_ _06100_ net389 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13167_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__inv_2
XANTENNA__12442__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ _05236_ _06031_ _05194_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ net325 net2161 net586 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13098_ _07072_ net227 _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12049_ net306 net2421 net531 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10305__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07590_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] _03450_ vssd1 vssd1 vccd1
+ vccd1 _03481_ sky130_fd_sc_hd__or2_1
X_15808_ clknet_leaf_8_wb_clk_i _02259_ _00766_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_16788_ net1342 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15739_ clknet_leaf_119_wb_clk_i _02190_ _00697_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16464__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14893__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09260_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\] net852 net848 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a22o_1
XANTENNA__08891__A team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08211_ _04089_ _04090_ _04073_ _04076_ _04079_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_29_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09191_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] net724 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\]
+ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] team_02_WB.instance_to_wrap.top.a1.dataIn\[0\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09631__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ _03960_ _03930_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12352__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ net882 _04636_ _04639_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[21\] vssd1 vssd1 vccd1 vccd1
+ net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[27\] vssd1 vssd1 vccd1 vccd1
+ net1424 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[0\] vssd1 vssd1 vccd1 vccd1
+ net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03814_ _03815_ vssd1 vssd1
+ vccd1 vccd1 _03817_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold48 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[5\] vssd1 vssd1 vccd1 vccd1
+ net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[1\] vssd1 vssd1 vccd1 vccd1
+ net1457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07857_ _03746_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11492__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07788_ _03637_ _03643_ _03674_ _03641_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a22o_2
XFILLER_0_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09527_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[18\] net665 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09458_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] net685 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09870__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08409_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03417_ _04274_ vssd1 vssd1
+ vccd1 vccd1 _04276_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12527__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] net795 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13212__A team_02_WB.START_ADDR_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ net422 _06626_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08425__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10232__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13050__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ net421 _06536_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15981__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10302_ net376 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14070_ net1111 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
X_11282_ net414 _06418_ _06899_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08740__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12770__B _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11667__A team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _06776_ net226 _03042_ net888 _03040_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12262__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ _05887_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__and2_2
XFILLER_0_63_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10535__A2 _05174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1002 net1015 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
X_10164_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] net716 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\]
+ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_4
Xfanout1024 net1027 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_4
Xfanout1035 net1049 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_4
Xfanout1046 net1049 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1057 net1067 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_2
XFILLER_0_41_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10095_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\] net738 net666 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a22o_1
X_14972_ net1034 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
Xfanout1068 net1072 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_4
Xfanout1079 net1086 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XFILLER_0_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09153__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13923_ net1073 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_16711_ net1265 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XANTENNA__11606__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16642_ net1213 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ net1070 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _05633_ _05635_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16573_ clknet_leaf_88_wb_clk_i net1404 _01446_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13785_ net1060 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10997_ net450 _06414_ _06635_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a21o_1
X_15524_ clknet_leaf_53_wb_clk_i _01975_ _00482_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12736_ team_02_WB.instance_to_wrap.top.a1.state\[1\] _07359_ _07361_ _07356_ vssd1
+ vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09861__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15455_ clknet_leaf_27_wb_clk_i _01906_ _00413_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12437__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _06689_ _06765_ _07293_ _07294_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__or4b_1
XANTENNA__10746__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14406_ net1094 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
X_11618_ net286 net1817 net576 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
X_15386_ clknet_leaf_120_wb_clk_i _01837_ _00344_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12598_ net933 net996 _04345_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__or3b_1
XFILLER_0_53_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16800__1354 vssd1 vssd1 vccd1 vccd1 _16800__1354/HI net1354 sky130_fd_sc_hd__conb_1
X_14337_ net1103 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11549_ _06001_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__nand2_1
Xhold507 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold518 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold529 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ net1085 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16007_ clknet_leaf_14_wb_clk_i _02458_ _00965_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13219_ team_02_WB.START_ADDR_VAL_REG\[27\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net211 sky130_fd_sc_hd__a21o_1
XANTENNA__12172__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ net1108 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XANTENNA__09392__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08760_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[12\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[12\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_2
Xhold1218 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1229 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07711_ _03573_ _03579_ _03571_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__o21ai_1
X_08691_ net745 _04449_ _04466_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__and3_4
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07642_ _03523_ _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15854__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07573_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09312_ _04983_ _04985_ _04987_ _04989_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[24\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_53_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09852__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09243_ _04915_ _04917_ _04919_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__or4_4
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12347__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14128__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout329_A _07015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ _04848_ _04850_ _04852_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08125_ _03990_ _04006_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__xor2_4
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08056_ _03942_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or2_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08560__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout698_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12082__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09383__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput105 wbs_we_i vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout865_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] net886 vssd1 vssd1 vccd1
+ vccd1 _04643_ sky130_fd_sc_hd__nand2_1
XANTENNA__09135__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ _03798_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08889_ net1540 _04575_ net825 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__mux2_1
X_10920_ _06366_ _06374_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__nand2_1
XANTENNA__13219__A1 team_02_WB.START_ADDR_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10150__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ net387 _06487_ _06497_ net399 vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13570_ net1171 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09843__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10782_ _06430_ _06432_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[30\]
+ sky130_fd_sc_hd__or2_2
XFILLER_0_94_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ net1740 net312 net477 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
XANTENNA__10453__A1 _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12257__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15240_ clknet_leaf_18_wb_clk_i _01691_ _00198_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12452_ net291 net2577 net484 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ net429 _06997_ _06999_ net442 _07011_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[9\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15171_ clknet_leaf_45_wb_clk_i _01622_ _00129_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12383_ net323 net2614 net492 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07875__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14122_ net1014 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
X_11334_ _05482_ net432 _06947_ net438 _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__a221o_1
XANTENNA__08470__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14053_ net1087 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
X_11265_ _06283_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13004_ _07366_ _03028_ team_02_WB.instance_to_wrap.top.pc\[22\] net944 vssd1 vssd1
+ vccd1 vccd1 _01520_ sky130_fd_sc_hd__a2bb2o_1
X_10216_ _05865_ _05867_ _05869_ _05871_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__or4_1
XANTENNA__09374__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11196_ net435 _06820_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] net775 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09126__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14955_ net999 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
X_10078_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\] net775 net842 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ net1081 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
X_14886_ net1167 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XANTENNA__10141__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13837_ net1132 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
X_16625_ clknet_leaf_67_wb_clk_i _02859_ _01498_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15107__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12969__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16556_ clknet_leaf_37_wb_clk_i net1436 _01429_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13768_ net1096 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
XANTENNA__09834__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12719_ _04578_ _04579_ _04666_ _07345_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__and4bb_1
X_15507_ clknet_leaf_124_wb_clk_i _01958_ _00465_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12167__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16487_ clknet_leaf_84_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[22\] _01361_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ net1071 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15438_ clknet_leaf_33_wb_clk_i _01889_ _00396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15369_ clknet_leaf_29_wb_clk_i _01820_ _00327_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 team_02_WB.instance_to_wrap.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net1702
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold315 team_02_WB.instance_to_wrap.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net1713
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 net115 vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold337 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold348 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net749 _05592_ vssd1
+ vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__o21a_2
Xhold359 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 _04658_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09365__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] net734 net714 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout817 net820 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_6
Xfanout828 _03297_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_4
Xfanout839 _04676_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_8
X_08812_ net183 net951 net902 net1499 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
Xhold1004 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] net692 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a22o_1
Xhold1015 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1026 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09117__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ net1645 net958 net924 _04528_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
Xhold1037 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1059 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08674_ net745 _04446_ _04466_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__and3_4
XFILLER_0_36_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08876__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _03446_ _03477_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12866__A team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07556_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] _03444_ vssd1 vssd1 vccd1
+ vccd1 _03447_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08555__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12077__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] team_02_WB.instance_to_wrap.ramload\[18\]
+ net967 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] net856 net778 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13385__B1 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09157_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] net700 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08108_ _03959_ _03966_ _03964_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a21oi_1
X_09088_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] net786 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout982_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08039_ _03892_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand2_2
Xhold860 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net403 _06364_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__or2_1
Xhold893 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10001_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\] net712 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12540__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09108__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14740_ net1200 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11952_ net284 net1844 net536 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10903_ team_02_WB.instance_to_wrap.top.pc\[27\] _06343_ vssd1 vssd1 vccd1 vccd1
+ _06547_ sky130_fd_sc_hd__xnor2_1
X_14671_ net1043 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11883_ net319 net2258 net546 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16410_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[9\]
+ _01284_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ net1106 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ _06048_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__or2_1
XANTENNA__16525__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16341_ clknet_leaf_100_wb_clk_i _02774_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13553_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] _03387_
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] vssd1 vssd1 vccd1
+ vccd1 _03390_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10765_ net379 _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ net2217 net257 net478 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__mux2_1
X_16272_ clknet_leaf_97_wb_clk_i _02705_ _01224_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13484_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] _03132_ vssd1 vssd1 vccd1 vccd1
+ _03345_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10696_ _06319_ _06327_ _06347_ team_02_WB.instance_to_wrap.top.aluOut\[31\] net461
+ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__o32a_4
XFILLER_0_129_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15223_ clknet_leaf_120_wb_clk_i _01674_ _00181_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12435_ net242 net2707 net485 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09595__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ clknet_leaf_25_wb_clk_i _01605_ _00112_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12366_ net234 net2568 net499 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14105_ net1062 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ net908 _06278_ _06929_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ clknet_leaf_77_wb_clk_i _01536_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ net354 net2629 net507 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__mux2_1
X_14036_ net1053 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XANTENNA__09347__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _05399_ _06025_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__nor2_1
XANTENNA__08555__A0 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11179_ net442 _06787_ _06805_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[18\]
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_78_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16055__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15987_ clknet_leaf_125_wb_clk_i _02438_ _00945_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11066__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14938_ net1047 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XANTENNA__10114__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08858__B2 net1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14869_ net1186 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ clknet_leaf_69_wb_clk_i _02842_ _01481_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ net1755 net935 net918 _04261_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09060__A _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ clknet_leaf_0_wb_clk_i net1431 _01412_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__A _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09011_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] net777 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ _04683_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[8\] vssd1 vssd1 vccd1
+ vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[25\] vssd1 vssd1 vccd1
+ vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold123 team_02_WB.instance_to_wrap.top.pc\[1\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\] vssd1
+ vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 team_02_WB.instance_to_wrap.top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1 net1543
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _02603_ vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold167 team_02_WB.instance_to_wrap.top.pc\[6\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] net730 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a221o_1
Xhold178 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[10\] vssd1 vssd1 vccd1
+ vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout625 net627 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _04488_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_8
X_09844_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\] net824 net820 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a22o_1
Xfanout647 _04486_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_2
XANTENNA__12360__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1103_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__A2_N _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _04477_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_4
X_09775_ _05421_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[29\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[29\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_1
XANTENNA__08849__A1 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10105__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15422__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16548__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] _04439_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07608_ _03467_ _03468_ _03473_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__and3_1
X_08588_ net973 _04373_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07539_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ _03429_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15572__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11005__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10550_ _04972_ _04990_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16679__1233 vssd1 vssd1 vccd1 vccd1 _16679__1233/HI net1233 sky130_fd_sc_hd__conb_1
XFILLER_0_134_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12535__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10481_ _04601_ _04602_ _06130_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14316__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ net283 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\] net513 vssd1
+ vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__mux2_1
XANTENNA__09577__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ net325 net1806 net520 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11102_ net404 _06494_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net305 net2086 net526 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
Xhold690 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16078__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033_ _04629_ net743 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] net443
+ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__a221o_1
X_15910_ clknet_leaf_13_wb_clk_i _02361_ _00868_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12270__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14051__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15841_ clknet_leaf_130_wb_clk_i _02292_ _00799_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ clknet_leaf_63_wb_clk_i _02223_ _00730_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ team_02_WB.instance_to_wrap.top.pc\[25\] net943 _03009_ _03011_ vssd1 vssd1
+ vccd1 vccd1 _01523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11844__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14723_ net1042 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
X_11935_ net239 net2122 net537 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output113_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14654_ net1033 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
X_11866_ net360 net1858 net548 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10738__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13605_ net1073 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
X_10817_ _06461_ _06465_ net388 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__a21oi_1
X_14585_ net1061 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ net356 net1969 net559 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13536_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\]
+ _03376_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__and3_1
X_16324_ clknet_leaf_98_wb_clk_i _02757_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10748_ _06397_ _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12953__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16255_ clknet_leaf_93_wb_clk_i _02693_ _01212_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_109_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12445__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ net1176 _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__nor3_1
XANTENNA__10754__A _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10679_ team_02_WB.instance_to_wrap.top.pc\[8\] _06330_ vssd1 vssd1 vccd1 vccd1 _06331_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15206_ clknet_leaf_13_wb_clk_i _01657_ _00164_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09568__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12418_ net283 net2514 net488 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__mux2_1
X_16186_ clknet_leaf_63_wb_clk_i _02632_ _01144_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13398_ _03291_ _03401_ _03137_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__mux2_1
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput217 net217 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
X_15137_ clknet_leaf_0_wb_clk_i _01588_ _00095_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ net320 net2500 net498 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15068_ clknet_leaf_85_wb_clk_i _01519_ _00031_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ net1068 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12180__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _03749_ _03779_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__nor3_1
XANTENNA__15445__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14896__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\] net818 net802 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\]
+ _05217_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08894__A team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13285__C1 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__or2_1
X_09491_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\] net698 net686 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\]
+ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a221o_1
XANTENNA__07503__A1 team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ _04301_ net1586 net827 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__B _05174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08373_ _04235_ _04236_ _04243_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or3_1
XANTENNA__13052__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10810__A1 _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12355__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout311_A _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09559__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08767__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16220__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
XANTENNA_fanout680_A _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_2
XANTENNA_fanout778_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_2
XANTENNA__12090__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16501__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _06126_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout444 _06322_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_2
XANTENNA__10326__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 _06129_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
Xfanout466 _07225_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09192__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] net727 net663 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\]
+ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout477 _07224_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_6
Xfanout499 _07219_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] net817 net793 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\]
+ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08709_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04367_ _04426_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09689_ _05337_ _05355_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11720_ net283 net2725 net566 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ net267 net2007 net572 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
X_10602_ net928 _05679_ net590 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14370_ net1091 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09798__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11582_ net380 _06403_ _07172_ net392 vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13321_ _03209_ _03221_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__and2b_1
X_10533_ _05238_ _05318_ _06184_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12265__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ clknet_leaf_55_wb_clk_i _02491_ _00998_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13252_ team_02_WB.instance_to_wrap.ramload\[25\] net980 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[25\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input74_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ _06101_ _06116_ net403 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ net237 net2459 net512 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13183_ _03167_ _03168_ _03149_ _03163_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10395_ _04826_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__and2_1
XANTENNA__08979__A team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ net236 net1912 net588 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11609__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ net356 net2601 net531 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10317__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ net414 _06424_ _06651_ _06411_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__a31o_1
XANTENNA__10868__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08930__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15824_ clknet_leaf_39_wb_clk_i _02275_ _00782_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12967_ _02867_ _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__xnor2_1
X_15755_ clknet_leaf_15_wb_clk_i _02206_ _00713_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10749__A _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07497__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10096__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ net270 net1903 net540 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
X_14706_ net1033 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15686_ clknet_leaf_12_wb_clk_i _02137_ _00644_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12898_ _02928_ _02931_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14637_ net1164 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
X_11849_ net318 net2555 net550 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09789__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14568_ net1099 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08997__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__A2 team_02_WB.instance_to_wrap.top.aluOut\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16307_ clknet_leaf_80_wb_clk_i _02740_ _01250_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13519_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03366_
+ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and2_1
XANTENNA__12175__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14499_ net1023 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16238_ clknet_leaf_71_wb_clk_i _00008_ _01195_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08749__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ clknet_leaf_71_wb_clk_i _02615_ _01127_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07793__A team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08991_ net882 _04639_ _04651_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__and3_4
XFILLER_0_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11519__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ _03764_ _03817_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03756_ vssd1 vssd1 vccd1
+ vccd1 _03764_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16678__1232 vssd1 vssd1 vccd1 vccd1 _16678__1232/HI net1232 sky130_fd_sc_hd__conb_1
XANTENNA__08921__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] net680 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09543_ _05205_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nor2_8
XANTENNA_fanout261_A _06586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07488__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] net789 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold1007_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ net960 _04285_ _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1170_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _04229_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12085__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _04162_ _04164_ _04157_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_85_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15610__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout895_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10011__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ net412 _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15760__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout241 _03894_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_4
Xfanout252 _06521_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_2
XANTENNA__09704__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net266 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
Xfanout274 _06674_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout285 _06912_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 _06753_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_1
XANTENNA__11511__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ net1064 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12768__B _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12821_ _07389_ _07444_ _07387_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07479__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15540_ clknet_leaf_46_wb_clk_i _01991_ _00498_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12752_ _04972_ _06241_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10078__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ net240 net2643 net566 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15471_ clknet_leaf_35_wb_clk_i _01922_ _00429_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15140__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12683_ _06537_ _06603_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13016__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14422_ net1106 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11634_ net594 _04579_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__or3_4
XFILLER_0_33_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11578__A2 team_02_WB.instance_to_wrap.top.aluOut\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14353_ net1029 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_11565_ net423 _06822_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15290__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ net985 _03400_ _03207_ _03209_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10516_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__inv_2
XANTENNA__10250__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14284_ net1002 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
X_11496_ _06397_ _06400_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13235_ team_02_WB.instance_to_wrap.ramload\[8\] net982 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[8\]
+ sky130_fd_sc_hd__and2_1
X_16023_ clknet_leaf_116_wb_clk_i _02474_ _00981_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ _06096_ _06099_ net364 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10002__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09943__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ _02782_ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10378_ _05238_ _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ net321 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\] net589 vssd1
+ vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
X_13097_ net230 _03104_ _03105_ _07425_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09156__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12048_ net298 net2185 net528 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15807_ clknet_leaf_10_wb_clk_i _02258_ _00765_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16787_ net1341 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XANTENNA__10479__A _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ net1126 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XANTENNA__10069__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15738_ clknet_leaf_120_wb_clk_i _02189_ _00696_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15669_ clknet_leaf_115_wb_clk_i _02120_ _00627_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08891__B _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _04076_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09190_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] net653 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15633__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _04001_ _04002_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _03910_ _03926_ _03932_ _03933_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a22o_1
XANTENNA__10241__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09934__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08974_ _04645_ _04653_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[3\] vssd1 vssd1 vccd1 vccd1
+ net1414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07925_ _03814_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__or2_1
Xhold27 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[7\] vssd1 vssd1 vccd1 vccd1
+ net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[25\] vssd1 vssd1 vccd1 vccd1
+ net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[3\] vssd1 vssd1 vccd1 vccd1
+ net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout476_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _03710_ _03715_ _03719_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07787_ _03660_ _03671_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout643_A _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] net733 net706 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__a221o_1
XANTENNA__11257__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] net716 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout810_A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11712__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ net990 _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09388_ _05057_ _05059_ _05061_ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13212__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08339_ net1680 net938 net920 _04215_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XANTENNA__08425__A2 _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11350_ net402 _06961_ _06962_ net412 vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ net898 _05936_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11281_ net414 _06426_ _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12543__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09386__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ _07446_ _03041_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__xor2_1
X_10232_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] _04427_ net749 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11667__B team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 net1006 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_4
X_10163_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] net652 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1014 net1015 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09138__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 net1027 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_2
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_4
XANTENNA_input37_A wbm_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1049 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_4
X_14971_ net1048 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
X_10094_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net714 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a221o_1
Xfanout1058 net1066 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_4
Xfanout1069 net1072 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
X_16710_ net1264 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13922_ net1089 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16641_ net1212 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ net1055 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14994__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12804_ _07406_ _07425_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o21a_1
X_16572_ clknet_leaf_91_wb_clk_i net1409 _01445_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ net1057 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
X_10996_ net413 _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__and2_1
XANTENNA__15656__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09310__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15523_ clknet_leaf_42_wb_clk_i _01974_ _00481_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12735_ _07352_ _07355_ _07359_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11622__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ net417 _06850_ _06820_ _06801_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__o211a_1
X_15454_ clknet_leaf_5_wb_clk_i _01905_ _00412_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10746__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ net1087 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
X_11617_ net269 net1726 net576 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XANTENNA__13122__B net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15385_ clknet_leaf_117_wb_clk_i _01836_ _00343_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12597_ net234 net2174 net475 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10223__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16677__1231 vssd1 vssd1 vccd1 vccd1 _16677__1231/HI net1231 sky130_fd_sc_hd__conb_1
XFILLER_0_135_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11548_ _05976_ _06000_ _05934_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_29_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14336_ net1083 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold508 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ net1060 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
Xhold519 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12453__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11479_ _06103_ _06105_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__nand2_1
XANTENNA__10762__A _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16006_ clknet_leaf_13_wb_clk_i _02457_ _00964_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13218_ team_02_WB.START_ADDR_VAL_REG\[26\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net210 sky130_fd_sc_hd__a21o_1
XFILLER_0_106_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09916__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14198_ net1106 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XANTENNA__10481__B _04602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13149_ net896 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09129__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1208 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16431__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ _03596_ _03600_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__nor2_1
X_08690_ net746 _04443_ _04446_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__and3_4
XANTENNA_wire611_A _05071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _03491_ _03524_ _03529_ _03530_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__and4b_1
XFILLER_0_75_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _03457_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16581__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09301__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] net790 net879 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10937__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\] net711 net684 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\]
+ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] net818 net813 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\]
+ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08124_ _03990_ _04006_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__nand2_1
XANTENNA__10214__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11465__A2_N net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03932_ _03933_ vssd1 vssd1
+ vccd1 vccd1 _03943_ sky130_fd_sc_hd__and3_1
XANTENNA__12363__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1133_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09368__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08142__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15529__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08957_ net882 _04639_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout760_A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11707__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _03787_ _03793_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__xnor2_1
X_08888_ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] net940 _04328_ net990 _04574_
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09540__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ _03717_ _03718_ _03686_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10850_ net387 _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] net844 net836 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10781_ net441 _06349_ _06431_ net428 vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__a22o_1
XANTENNA__12538__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12520_ net2074 net310 net479 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ net283 net2283 net485 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ net434 _07005_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15170_ clknet_leaf_48_wb_clk_i _01621_ _00128_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12382_ net319 net2210 net495 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12781__B _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ net1012 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ _05484_ net455 net446 _05483_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__a22o_1
XANTENNA__12273__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14054__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09359__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ net1143 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
X_11264_ _06269_ _06281_ _06282_ _04416_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__a31o_1
XANTENNA__14989__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13003_ _06696_ net226 _03027_ net888 _03026_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__o221a_1
X_10215_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] net695 net659 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11195_ net409 _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10146_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\] net837 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] net855 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__a22o_1
X_14954_ net1009 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09531__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ net1029 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
X_14885_ net1165 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
X_16624_ clknet_leaf_60_wb_clk_i _02858_ _01497_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13836_ net1005 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16555_ clknet_leaf_7_wb_clk_i net1434 _01428_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10979_ net264 net2677 net583 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
X_13767_ net1152 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XANTENNA__12448__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13091__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15506_ clknet_leaf_25_wb_clk_i _01957_ _00464_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12718_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] net974 team_02_WB.instance_to_wrap.top.a1.instruction\[11\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1 vccd1 vccd1 _07345_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ clknet_leaf_85_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[21\] _01360_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08227__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13698_ net1092 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15437_ clknet_leaf_21_wb_clk_i _01888_ _00395_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12649_ _04992_ _05032_ _05074_ _05114_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15368_ clknet_leaf_110_wb_clk_i _01819_ _00326_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09062__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12183__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14319_ net1123 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold305 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold316 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ clknet_leaf_40_wb_clk_i _01750_ _00257_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold327 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 team_02_WB.instance_to_wrap.top.a1.row1\[12\] vssd1 vssd1 vccd1 vccd1 net1736
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09860_ _05503_ _05521_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__nor2_2
Xfanout807 _04658_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
Xfanout818 net820 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
Xfanout829 net832 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15821__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ net184 net951 net902 net1490 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
XANTENNA__09770__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] net730 net666 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\]
+ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a221o_1
Xhold1005 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1027 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[21\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[21\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_2
Xhold1038 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1049 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ net748 _04442_ _04466_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__and3_1
XANTENNA__15971__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07624_ _03478_ _03479_ _03506_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07555_ _03444_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
XANTENNA__12358__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1083_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07486_ net2732 team_02_WB.instance_to_wrap.ramload\[19\] net967 vssd1 vssd1 vccd1
+ vccd1 _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] net836 net758 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09589__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] net715 net662 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\]
+ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09053__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08107_ _03959_ _03964_ net225 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\] net858 net834 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a22o_1
XANTENNA__16504__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12093__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08800__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08038_ _03882_ _03886_ net241 vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold850 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold872 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold894 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\] net716 net685 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a22o_1
XANTENNA__09761__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09989_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] net855 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16676__1230 vssd1 vssd1 vccd1 vccd1 _16676__1230/HI net1230 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11951_ net270 net2137 net536 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10902_ net441 _06523_ _06543_ _06546_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[27\]
+ sky130_fd_sc_hd__a211o_2
X_11882_ net317 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\] net545 vssd1
+ vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
X_14670_ net1033 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08746__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13621_ net1114 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
X_10833_ _04826_ _06047_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16340_ clknet_leaf_100_wb_clk_i _02773_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13552_ net1603 _03387_ _03389_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10764_ _04625_ net371 _06370_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09292__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12503_ net1769 net252 net478 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13483_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ _03132_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _03344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16271_ clknet_leaf_93_wb_clk_i _02704_ _01223_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net912 _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nor2_1
XANTENNA__11900__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12434_ net237 net1911 net484 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__mux2_1
X_15222_ clknet_leaf_110_wb_clk_i _01673_ _00180_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09044__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15153_ clknet_leaf_17_wb_clk_i _01604_ _00111_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12365_ net361 net2291 net497 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__mux2_1
XANTENNA__13400__B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14104_ net1063 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_11316_ net913 _06931_ _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1
+ vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__a2bb2o_1
X_15084_ clknet_leaf_77_wb_clk_i _01535_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15844__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ net343 net2354 net504 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14035_ net1148 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11247_ net427 _06867_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09752__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__A _05257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net428 _06788_ _06796_ net451 _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15994__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10129_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\] net815 net766 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ clknet_leaf_25_wb_clk_i _02437_ _00944_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09504__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14937_ net1043 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XANTENNA__08858__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15224__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14868_ net1186 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
X_16607_ clknet_leaf_83_wb_clk_i _02841_ _01480_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ net1047 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12178__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13064__B1 _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ net1198 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16538_ clknet_leaf_129_wb_clk_i net1458 _01411_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09060__B _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09283__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15374__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13798__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ clknet_leaf_99_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[4\] _01343_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09010_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\] net878 _04693_ _04694_
+ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09035__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold102 _02587_ vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold113 _02604_ vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__B net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10050__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold124 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[0\] vssd1 vssd1 vccd1
+ vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09991__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[13\] vssd1 vssd1 vccd1
+ vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold146 team_02_WB.instance_to_wrap.top.pc\[28\] vssd1 vssd1 vccd1 vccd1 net1544
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 team_02_WB.instance_to_wrap.top.a1.data\[6\] vssd1 vssd1 vccd1 vccd1 net1555
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold168 net114 vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\] net726 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__a22o_1
Xhold179 _02589_ vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout615 _04425_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_4
Xfanout626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_6
XANTENNA__09743__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] net788 net764 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a221o_1
Xfanout637 _04488_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_4
Xfanout648 net651 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_6
Xfanout659 _04481_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA_fanout389_A _05908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[13\] net592 vssd1
+ vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_119_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08725_ net1643 net955 net924 _04519_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08849__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _07197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ net746 _04443_ _04449_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07607_ _03483_ _03488_ _03495_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08587_ net979 _04369_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and2_1
XANTENNA__12088__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15717__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07538_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] team_02_WB.instance_to_wrap.top.a1.dataIn\[26\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__or4_1
XFILLER_0_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07469_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _03409_
+ sky130_fd_sc_hd__inv_2
XANTENNA__08482__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11720__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09208_ _04878_ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10480_ net580 net448 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09026__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] net879 net754 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\]
+ _04805_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08785__B2 _04549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ net319 net2464 net523 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XANTENNA__09982__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11101_ net398 _06490_ _06731_ net411 vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12081_ net296 net1829 net524 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
XANTENNA__12551__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _06341_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__or2_1
XANTENNA__11541__A0 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A1 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15840_ clknet_leaf_12_wb_clk_i _02291_ _00798_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ clknet_leaf_105_wb_clk_i _02222_ _00729_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__inv_2
XANTENNA__12787__A _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14722_ net1008 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
X_11934_ _07192_ _07199_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13046__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ net1007 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
XANTENNA__16409__D team_02_WB.instance_to_wrap.top.ru.dmmload_co\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ net353 net1988 net548 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13604_ net1100 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10816_ net375 _06419_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14584_ net1062 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11796_ net344 net2215 net557 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__mux2_1
XANTENNA__09265__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16323_ clknet_leaf_98_wb_clk_i _02756_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ _03377_ _03378_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nor2_1
X_10747_ _05722_ net369 vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__nand2_1
XANTENNA__11630__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16254_ clknet_leaf_98_wb_clk_i _02692_ _01211_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_13466_ net1547 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03331_ vssd1
+ vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__and3_1
X_10678_ team_02_WB.instance_to_wrap.top.pc\[7\] team_02_WB.instance_to_wrap.top.pc\[6\]
+ _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15205_ clknet_leaf_125_wb_clk_i _01656_ _00163_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12417_ net267 net2576 net488 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__mux2_1
X_16185_ clknet_leaf_66_wb_clk_i _02631_ _01143_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
X_13397_ net1724 net896 _03295_ net993 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__o211a_1
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XANTENNA__10032__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput218 net218 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_15136_ clknet_leaf_7_wb_clk_i _01587_ _00094_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12348_ net317 net2731 net497 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12461__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net289 net2081 net504 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__mux2_1
X_15067_ clknet_leaf_84_wb_clk_i _01518_ _00030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14242__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ net1091 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15969_ clknet_leaf_2_wb_clk_i _02420_ _00927_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__nor2_4
XANTENNA__08894__B team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09490_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] net723 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08441_ net960 _04299_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08372_ net1699 net935 net918 _04245_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XANTENNA__09256__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11540__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10271__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout304_A _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1046_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__B2 _04540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14152__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
XANTENNA__16515__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 _05817_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09716__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_2
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_A _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout445 net447 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13991__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 _04505_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout467 _07225_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_4
X_09826_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] net723 net667 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 _07224_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 net491 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_6
XFILLER_0_57_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout840_A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] net857 net777 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11715__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08708_ net928 net462 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nor2_1
X_09688_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13028__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ _04364_ _04368_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_132_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11650_ net324 net2582 net572 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XANTENNA__09247__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ net928 _05545_ net590 vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11581_ _04502_ net369 vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nand2_1
XANTENNA__12546__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13231__A team_02_WB.instance_to_wrap.ramload\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10262__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13320_ _03218_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__nor2_4
XFILLER_0_49_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10532_ _05277_ _06028_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nor2_2
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07695__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16045__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13251_ net1692 net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[24\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10463_ _06107_ _06115_ net390 vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _04428_ _04579_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__or3b_4
XFILLER_0_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09955__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ _03146_ _02780_ _03166_ _02785_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a31o_1
XANTENNA_input67_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10394_ _04911_ _06046_ _04867_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ net360 net1868 net586 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XANTENNA__12281__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09707__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net342 net2107 net528 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__mux2_1
XANTENNA__08060__A team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ _06424_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout990 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1
+ net990 sky130_fd_sc_hd__buf_2
X_15823_ clknet_leaf_34_wb_clk_i _02274_ _00781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11625__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15754_ clknet_leaf_44_wb_clk_i _02205_ _00712_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09486__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10749__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ net1186 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _06856_ net2140 net540 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15685_ clknet_leaf_125_wb_clk_i _02136_ _00643_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08694__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ team_02_WB.instance_to_wrap.top.pc\[2\] _05936_ _02930_ vssd1 vssd1 vccd1
+ vccd1 _02931_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ net1166 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ net303 net2499 net551 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XANTENNA__09238__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ net1153 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
XANTENNA__12456__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11779_ net290 net2327 net556 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16306_ clknet_leaf_80_wb_clk_i _02739_ _01249_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13518_ _03366_ _03367_ net885 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__and3b_1
X_14498_ net1090 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16237_ clknet_leaf_70_wb_clk_i _00007_ _01194_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] _03321_ net1671 vssd1 vssd1
+ vccd1 vccd1 _03324_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10005__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15412__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09946__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16168_ clknet_leaf_71_wb_clk_i _02614_ _01126_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09410__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15119_ clknet_leaf_35_wb_clk_i _01570_ _00077_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12191__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16099_ clknet_leaf_70_wb_clk_i _02545_ _01057_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08990_ _04633_ _04636_ _04639_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and3_1
XANTENNA__07972__A2 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _03817_ _03818_ net262 vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a21boi_1
XANTENNA__15562__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07872_ _03760_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire906_A _04552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] net712 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[16\]
+ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09542_ _05207_ _05209_ _05211_ _05213_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__or4_2
XFILLER_0_56_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09477__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ _05141_ _05143_ _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08685__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08424_ team_02_WB.instance_to_wrap.top.a1.row1\[19\] net827 vssd1 vssd1 vccd1 vccd1
+ _04289_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _04225_ _04228_ _04220_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout421_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout519_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10244__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _04165_ _03425_ net937 net2711 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15092__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09937__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout790_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10547__A1 _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09401__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15905__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16512__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xfanout253 _06521_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_1
XFILLER_0_22_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout264 net266 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 _06912_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_1
Xfanout297 _06753_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\] net867 net851 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ _07388_ _07443_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10569__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12751_ _04932_ _06237_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11702_ net594 _04578_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__or3_4
X_15470_ clknet_leaf_39_wb_clk_i _01921_ _00428_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08754__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12682_ _04625_ net448 _06423_ _06464_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__or4_1
XANTENNA__12784__B _05797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14421_ net1121 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04428_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12276__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10235__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14352_ net1017 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
Xwire610 _05112_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08055__A team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11564_ net398 _07003_ _07156_ net411 vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09640__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ net986 net987 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__nand2b_1
X_10515_ _05678_ _05700_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__a21o_1
X_11495_ net346 net2524 net584 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14283_ net1014 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16022_ clknet_leaf_112_wb_clk_i _02473_ _00980_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ team_02_WB.instance_to_wrap.ramload\[7\] net982 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[7\]
+ sky130_fd_sc_hd__and2_1
X_10446_ _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13165_ _03153_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__inv_2
X_10377_ _06027_ _06029_ _05276_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__o21a_1
X_12116_ net316 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\] net587 vssd1
+ vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
X_13096_ _07407_ _07422_ _07424_ net890 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_40_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12047_ net287 net2319 net528 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15806_ clknet_leaf_4_wb_clk_i _02257_ _00764_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ net1340 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
X_13998_ net1115 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15737_ clknet_leaf_108_wb_clk_i _02188_ _00695_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12949_ net229 _02980_ net226 _06436_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08667__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15668_ clknet_leaf_49_wb_clk_i _02119_ _00626_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14619_ net1193 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12186__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ clknet_leaf_33_wb_clk_i _02050_ _00557_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08140_ _03988_ _04011_ _04014_ _04024_ _04009_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09092__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10777__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ _03940_ _03950_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21bo_1
XANTENNA__15928__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09919__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11726__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08973_ net882 _04636_ _04644_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and3_4
XFILLER_0_80_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold17 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[19\] vssd1 vssd1 vccd1 vccd1
+ net1415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07924_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03790_ _03791_ vssd1 vssd1
+ vccd1 vccd1 _03815_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold28 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[4\] vssd1 vssd1 vccd1 vccd1
+ net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[13\] vssd1 vssd1 vccd1 vccd1
+ net1437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09524__A _05175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07855_ _03710_ _03714_ _03719_ _03711_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a31o_1
XANTENNA__15308__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ _03675_ _03676_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] net694 net662 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout636_A _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15458__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\] net668 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\]
+ _05129_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08407_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] team_02_WB.instance_to_wrap.top.a1.halfData\[2\]
+ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__12096__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09387_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] net789 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\]
+ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10217__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08338_ _04199_ _04200_ _04209_ _04211_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__a41o_2
XANTENNA__09083__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08269_ _04122_ _04147_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__xor2_2
XANTENNA__08830__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[1\] vssd1 vssd1 vccd1
+ vccd1 _05954_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net412 _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__nand2_1
X_10231_ net462 _05841_ _05886_ net456 net740 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11667__C _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] net730 net709 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\]
+ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 net1067 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1026 net1027 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_4
X_14970_ net1043 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
Xfanout1037 net1049 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_2
X_10093_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\] net650 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a22o_1
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14340__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1066 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_2
X_13921_ net1144 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ net1211 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_13852_ net1097 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12803_ _07405_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16571_ clknet_leaf_89_wb_clk_i net1399 _01444_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13783_ net1115 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
X_10995_ net402 _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11903__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15522_ clknet_leaf_49_wb_clk_i _01973_ _00480_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12734_ _07352_ _07354_ _07360_ team_02_WB.instance_to_wrap.top.a1.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09861__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15453_ clknet_leaf_113_wb_clk_i _01904_ _00411_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12665_ _06716_ _06740_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10208__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14404_ net1093 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11616_ _06856_ net1710 net576 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XANTENNA__09074__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15384_ clknet_leaf_126_wb_clk_i _01835_ _00342_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09613__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ net360 net2628 net472 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14335_ net1118 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11547_ net422 _06797_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold509 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14266_ net1059 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08513__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11478_ net442 _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ clknet_leaf_127_wb_clk_i _02456_ _00963_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13217_ team_02_WB.START_ADDR_VAL_REG\[25\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net209 sky130_fd_sc_hd__a21o_1
X_10429_ _04972_ net373 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__nand2_1
X_14197_ net1120 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13148_ _03133_ _03138_ _03139_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_57_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13079_ net230 _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1209 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11593__B _04602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__A2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07640_ _03491_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15600__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07571_ _03438_ _03456_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1
+ vccd1 vccd1 _03462_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16769_ net1323 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] net863 net806 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__a22o_1
XANTENNA__11813__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09852__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\] net674 net653 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15750__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13397__C1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09172_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] net854 net850 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a22o_1
XANTENNA__09065__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _04005_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08812__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16106__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ _03932_ _03933_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1
+ vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08142__B team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15130__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_A _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08956_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07907_ _03783_ _03792_ _03797_ _03778_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12675__A1 _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net990 net916 _04321_ _04273_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07838_ _03727_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10150__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07769_ _03650_ _03653_ _03657_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_6_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11723__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09508_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\] net840 net756 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\]
+ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _04744_ _06213_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__xor2_1
XANTENNA__09843__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09439_ net897 net610 _04630_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__C1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09056__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net267 net2383 net484 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11401_ net449 _07006_ _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08803__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ net316 net2528 net493 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XANTENNA__12554__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__A2 _07005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14120_ net1096 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11332_ net423 _06495_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ net1068 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
X_11263_ net442 _06870_ _06883_ _06868_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[15\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13002_ _07380_ _07450_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10214_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\] net631 net623 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a22o_1
X_11194_ net400 _06604_ _06818_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10145_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\] net803 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07790__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15623__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10076_ _05729_ _05731_ _05733_ _05735_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__or4_1
XANTENNA__11469__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14953_ net1010 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13904_ net1017 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
X_14884_ net1162 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10141__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ clknet_leaf_65_wb_clk_i _02857_ _01496_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_13835_ net1014 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XANTENNA__15773__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12969__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ clknet_leaf_7_wb_clk_i net1433 _01427_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09295__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ net1139 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ _06615_ _06616_ _06617_ team_02_WB.instance_to_wrap.top.aluOut\[25\] net460
+ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__o32a_2
XFILLER_0_58_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09834__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15505_ clknet_leaf_16_wb_clk_i _01956_ _00463_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12717_ net988 _07343_ _07344_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16485_ clknet_leaf_86_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[20\] _01359_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13697_ net1144 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15436_ clknet_leaf_22_wb_clk_i _01887_ _00394_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09047__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12648_ _05155_ _05194_ _05237_ _05276_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15367_ clknet_leaf_114_wb_clk_i _01818_ _00325_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ net315 net2463 net474 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14318_ net1115 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
XANTENNA__10601__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ clknet_leaf_49_wb_clk_i _01749_ _00256_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold317 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold328 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold339 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net1024 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout808 _04658_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout819 net820 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11808__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ net154 net951 net902 net1576 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
X_16769__1323 vssd1 vssd1 vccd1 vccd1 _16769__1323/HI net1323 sky130_fd_sc_hd__conb_1
X_09790_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] net722 net708 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1006 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net1634 net956 net925 _04527_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
Xhold1028 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1039 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08672_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\] net693 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07533__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _03479_ _03506_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07554_ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] _03435_ _03437_ vssd1 vssd1
+ vccd1 vccd1 _03445_ sky130_fd_sc_hd__and3_1
XANTENNA__09286__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07485_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] net2554 net966 vssd1
+ vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16725__1279 vssd1 vssd1 vccd1 vccd1 _16725__1279/HI net1279 sky130_fd_sc_hd__conb_1
X_09224_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] net823 net818 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\]
+ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12882__B _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12374__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\] net642 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout501_A _07218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10199__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08106_ _03971_ _03975_ _03982_ _03985_ _03991_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__o311a_1
X_09086_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\] net863 net802 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ _04766_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08037_ _03920_ _03924_ _03922_ _03918_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__and4b_1
XFILLER_0_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold840 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold851 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold862 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15646__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap581 _04591_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_1
Xhold873 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold895 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11718__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16520__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09988_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\] net880 _05647_ _05649_
+ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08939_ _04614_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__nor2_4
XANTENNA__15796__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11950_ _06856_ net1784 net536 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10901_ net427 _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ net305 net2513 net546 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XANTENNA__12549__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10858__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ net1038 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10832_ net248 net2609 net582 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09277__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09816__A2 _05480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] _03387_
+ net884 vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10763_ _06412_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12502_ net2689 net249 net478 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XANTENNA__10831__B1 team_02_WB.instance_to_wrap.top.aluOut\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09029__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16270_ clknet_leaf_79_wb_clk_i _02703_ _01222_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input97_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ _03137_ _03309_ _03343_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__and3_1
XANTENNA__08762__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10694_ team_02_WB.instance_to_wrap.top.pc\[31\] _06345_ vssd1 vssd1 vccd1 vccd1
+ _06346_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15176__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15221_ clknet_leaf_115_wb_clk_i _01672_ _00179_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ _04576_ _07190_ _07199_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__or3_4
XFILLER_0_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10593__A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12284__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16421__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ clknet_leaf_39_wb_clk_i _01603_ _00110_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12364_ net351 net2466 net496 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ net1108 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11315_ _06334_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__or2_1
X_15083_ clknet_leaf_77_wb_clk_i _01534_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ net348 net1797 net505 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14034_ net1079 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XANTENNA__09201__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246_ _06151_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11628__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _05238_ net453 _06800_ _06802_ _06803_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__a2111o_1
X_10128_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\] net822 net842 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22o_1
X_15985_ clknet_leaf_19_wb_clk_i _02436_ _00943_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10059_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] net726 net670 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a22o_1
X_14936_ net1002 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12459__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ net1171 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10768__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16606_ clknet_leaf_67_wb_clk_i _02840_ _01479_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_13818_ net1058 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09268__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14798_ net1198 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16537_ clknet_leaf_129_wb_clk_i net1449 _01410_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13749_ net1118 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XANTENNA__15519__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ clknet_leaf_81_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[3\] _01342_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11599__A team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15419_ clknet_leaf_105_wb_clk_i _01870_ _00377_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12194__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16399_ clknet_leaf_83_wb_clk_i team_02_WB.instance_to_wrap.top.ru.r1.nxt_dmmWen
+ _01273_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmWen sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15669__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[7\] vssd1 vssd1 vccd1
+ vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold114 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[19\] vssd1 vssd1 vccd1
+ vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08794__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 _02579_ vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold136 _02592_ vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14703__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold147 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[11\] vssd1 vssd1 vccd1
+ vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold158 team_02_WB.instance_to_wrap.top.a1.data\[3\] vssd1 vssd1 vccd1 vccd1 net1556
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\] net722 net666 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\]
+ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold169 team_02_WB.START_ADDR_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout616 net619 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_8
X_09842_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] net867 net848 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a22o_1
Xfanout627 _04493_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_4
Xfanout638 _04488_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout649 net651 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_4
XANTENNA__08420__B _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _05430_ _05439_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[13\]
+ sky130_fd_sc_hd__or2_4
XFILLER_0_77_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout284_A _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[30\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[30\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10105__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08655_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\] net738 net734 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\]
+ _04451_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a221o_1
XANTENNA__12369__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1193_A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout549_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07606_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03496_ vssd1 vssd1 vccd1
+ vccd1 _03497_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13054__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09259__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ net978 _04369_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03426_ vssd1 vssd1 vccd1
+ vccd1 _03428_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout716_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07468_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _04880_ _04882_ _04884_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__or4_2
XANTENNA__16515__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] net810 net798 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__a221o_1
XANTENNA__16594__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08785__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09069_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\] net733 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ net403 _06485_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__or2_1
X_12080_ net289 net2300 net524 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
Xhold670 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold681 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13229__A team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11031_ team_02_WB.instance_to_wrap.top.pc\[23\] _06340_ vssd1 vssd1 vccd1 vccd1
+ _06667_ sky130_fd_sc_hd__nor2_1
XANTENNA__11541__A1 _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15770_ clknet_leaf_120_wb_clk_i _02221_ _00728_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ net989 net911 _04437_ _06614_ net943 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12787__B _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input12_A wbm_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ net1040 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ net235 net2453 net541 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12279__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ net1001 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11864_ net354 net2455 net551 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13603_ net1073 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XANTENNA__11057__B1 _06688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ net413 net396 _06462_ _06414_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a31o_1
X_14583_ net1119 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ net346 net1926 net557 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11911__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16322_ clknet_leaf_97_wb_clk_i _02755_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13534_ net2724 _03376_ net885 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__o21ai_1
X_10746_ _05768_ net375 vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15811__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16768__1322 vssd1 vssd1 vccd1 vccd1 _16768__1322/HI net1322 sky130_fd_sc_hd__conb_1
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09670__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16253_ clknet_leaf_92_wb_clk_i _02691_ _01210_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03331_ net1547 vssd1
+ vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ team_02_WB.instance_to_wrap.top.pc\[5\] _06328_ vssd1 vssd1 vccd1 vccd1 _06329_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_129_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ clknet_leaf_55_wb_clk_i _01655_ _00162_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net323 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\] net488 vssd1
+ vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16184_ clknet_leaf_71_wb_clk_i _02630_ _01142_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09422__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13396_ team_02_WB.instance_to_wrap.top.a1.row1\[101\] _03285_ _03293_ _03294_ vssd1
+ vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XANTENNA__09973__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ clknet_leaf_24_wb_clk_i _01586_ _00093_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12347_ net305 net2141 net498 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput219 net219 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ clknet_leaf_84_wb_clk_i _01517_ _00029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12278_ net279 net1783 net504 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14017_ net1101 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
X_11229_ _06580_ _06851_ _06630_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13063__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724__1278 vssd1 vssd1 vccd1 vccd1 _16724__1278/HI net1278 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09489__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ clknet_leaf_10_wb_clk_i _02419_ _00926_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14919_ net1166 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XANTENNA__12189__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15341__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15899_ clknet_leaf_118_wb_clk_i _02350_ _00857_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16467__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08440_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[7\] net917 vssd1 vssd1 vccd1
+ vccd1 _04300_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08700__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08371_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15491__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09661__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11341__A2_N net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09413__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1039_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout402 _05862_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_2
Xfanout413 net415 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 _05816_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11523__A1 _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 _06121_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10326__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
X_09825_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] net703 _05489_ vssd1
+ vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a21o_1
XANTENNA_input4_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 _06326_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09192__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 net471 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout479 _07224_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09756_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\] net781 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\]
+ _05422_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__a221o_1
XANTENNA__07481__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ net976 net615 _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12099__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[15\] net592 vssd1
+ vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout833_A _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13028__A1 team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08638_ _04388_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15834__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08569_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] team_02_WB.instance_to_wrap.top.a1.instruction\[2\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[1\] team_02_WB.instance_to_wrap.top.a1.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__or4bb_2
XANTENNA__11731__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10600_ net928 _05545_ net590 vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_119_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11580_ _04600_ _04701_ _06128_ _06216_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09652__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ _05195_ _05196_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15984__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16823__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ net1730 net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[23\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ _06110_ _06114_ net365 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09404__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04429_ vssd1 vssd1 vccd1 vccd1
+ _07214_ sky130_fd_sc_hd__o31ai_2
XANTENNA__12562__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13181_ _03146_ _02780_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14343__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10871__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ _04913_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_1
XANTENNA__15214__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12132_ net352 net2236 net586 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12063_ net347 net2423 net530 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10317__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ net396 _06650_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15364__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11906__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15822_ clknet_leaf_42_wb_clk_i _02273_ _00780_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout991 _03414_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15753_ clknet_leaf_32_wb_clk_i _02204_ _00711_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12965_ _06547_ net226 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14704_ net1193 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
X_11916_ net319 net2324 net543 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ clknet_leaf_19_wb_clk_i _02135_ _00642_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ team_02_WB.instance_to_wrap.top.pc\[1\] _04510_ _02929_ vssd1 vssd1 vccd1
+ vccd1 _02930_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ net1162 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11847_ net297 net1913 net548 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11641__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ net1140 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XANTENNA__09643__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11778_ net282 net1937 net556 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13517_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03367_ sky130_fd_sc_hd__a21o_1
XANTENNA__08997__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16305_ clknet_leaf_80_wb_clk_i _02738_ _01248_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ net382 _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11450__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14497_ net1144 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16236_ clknet_leaf_70_wb_clk_i _02677_ _01193_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.busy_o
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13448_ net2326 _03321_ _03323_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16167_ clknet_leaf_72_wb_clk_i _02613_ _01125_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12472__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ clknet_leaf_33_wb_clk_i _01569_ _00076_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16098_ clknet_leaf_80_wb_clk_i _02544_ _01056_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15707__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03827_ _03828_ _03829_ vssd1
+ vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15049_ clknet_leaf_91_wb_clk_i _01500_ net995 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10308__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07871_ _03731_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11816__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] net660 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__a22o_1
XANTENNA__08921__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15857__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\] net684 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\]
+ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09472_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] net853 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ _05136_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ team_02_WB.instance_to_wrap.top.a1.data\[11\] net915 _04287_ vssd1 vssd1
+ vccd1 vccd1 _04288_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout247_A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _04220_ _04225_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__and3_1
XANTENNA__08437__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09634__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11441__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ _04157_ _04162_ _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15237__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12890__B _05797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13194__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout783_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout232 _07330_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout243 net245 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net257 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 net278 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
X_16767__1321 vssd1 vssd1 vccd1 vccd1 _16767__1321/HI net1321 sky130_fd_sc_hd__conb_1
XANTENNA__11726__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08912__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] net807 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a22o_1
Xfanout287 net290 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout298 _06753_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_1
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\] net720 net672 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ _05405_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12750_ _04932_ _06237_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09873__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] _04428_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__or3b_4
XFILLER_0_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16012__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ _07308_ _06921_ _06900_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__or3b_1
XANTENNA__14338__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14420_ net1051 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ net235 net2331 net577 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ net1124 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ net390 _07081_ _07154_ _07155_ net404 vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__a221o_1
Xwire611 _05071_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_2
X_16723__1277 vssd1 vssd1 vccd1 vccd1 _16723__1277/HI net1277 sky130_fd_sc_hd__conb_1
XFILLER_0_110_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ net985 _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nor2_1
XANTENNA__16162__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10514_ _05703_ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08770__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14282_ net1031 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[5\] _07093_ vssd1 vssd1 vccd1
+ vccd1 _07094_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16021_ clknet_leaf_116_wb_clk_i _02472_ _00979_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ net2226 net984 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[6\]
+ sky130_fd_sc_hd__and2_1
X_10445_ _05633_ net372 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nand2_1
XANTENNA__12292__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13164_ net992 _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ _05316_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output166_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12115_ net306 net2558 net589 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux2_1
X_13095_ _02923_ _02936_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09156__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ net279 net2587 net528 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XANTENNA__11636__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15805_ clknet_leaf_116_wb_clk_i _02256_ _00763_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ net1134 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_16785_ net1339 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08116__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12948_ _07367_ _07368_ _02871_ net888 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15736_ clknet_leaf_121_wb_clk_i _02187_ _00694_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09864__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12467__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ clknet_leaf_126_wb_clk_i _02118_ _00625_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12879_ team_02_WB.instance_to_wrap.top.pc\[11\] _05548_ vssd1 vssd1 vccd1 vccd1
+ _02913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12694__C _07321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14618_ net1193 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15598_ clknet_leaf_42_wb_clk_i _02049_ _00556_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14549_ net1119 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10777__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08070_ _03920_ _03955_ _03956_ _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__and4b_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16219_ clknet_leaf_38_wb_clk_i _02664_ _01176_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _04649_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__nor2_4
XFILLER_0_53_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14711__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07923_ _03790_ _03791_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1
+ vccd1 vccd1 _03814_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09147__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[14\] vssd1 vssd1 vccd1 vccd1
+ net1416 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold29 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[4\] vssd1 vssd1 vccd1 vccd1
+ net1427 sky130_fd_sc_hd__dlygate4sd3_1
X_07854_ _03710_ _03719_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09524__B _05193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16035__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _03634_ _03663_ _03665_ _03628_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout364_A _05956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13100__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _05175_ _05193_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__B _05725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09455_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] net728 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a22o_1
XANTENNA__10686__A team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12377__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09386_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] net785 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13997__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08337_ _04195_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ _04146_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout998_A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _04066_ _04068_ _04072_ _04081_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10230_ net974 _04425_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a21o_1
XANTENNA__09386__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10161_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\] net690 net650 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09138__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1019 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_4
Xfanout1027 net1032 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_4
X_10092_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\] net693 net673 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a221o_1
Xfanout1049 net1067 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
X_13920_ net1082 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XANTENNA__10153__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__C1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13851_ net1046 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _05678_ _05681_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__nor2_1
X_13782_ net1109 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
X_16570_ clknet_leaf_99_wb_clk_i net1425 _01443_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09846__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15402__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _06504_ _06632_ net385 vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__mux2_1
XANTENNA__16528__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__inv_2
X_15521_ clknet_leaf_2_wb_clk_i _01972_ _00479_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12287__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15452_ clknet_leaf_61_wb_clk_i _01903_ _00410_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12664_ _07158_ _07177_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ net1068 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ net319 net1759 net578 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15383_ clknet_leaf_119_wb_clk_i _01834_ _00341_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ net351 net2458 net472 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ net1023 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XANTENNA__13700__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11546_ net423 _06795_ _07140_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__a21o_1
XANTENNA__08821__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14265_ net1065 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11477_ _06012_ _07077_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16004_ clknet_leaf_18_wb_clk_i _02455_ _00962_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13216_ team_02_WB.START_ADDR_VAL_REG\[24\] _04356_ vssd1 vssd1 vccd1 vccd1 net208
+ sky130_fd_sc_hd__and2_1
XFILLER_0_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ _04932_ net371 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__nand2_1
X_14196_ net1038 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__and4bb_1
X_10359_ _05837_ _06008_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09129__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13078_ _02939_ _02941_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__xor2_1
XANTENNA__16058__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net339 net2049 net469 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08888__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10144__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07570_ _03432_ _03440_ _03454_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ net1322 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09301__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15719_ clknet_leaf_16_wb_clk_i _02170_ _00677_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12197__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16699_ net1253 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09240_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] net662 _04918_ vssd1
+ vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08407__C team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\] net858 net794 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\]
+ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ _03985_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__xnor2_2
X_16766__1320 vssd1 vssd1 vccd1 vccd1 _16766__1320/HI net1320 sky130_fd_sc_hd__conb_1
XFILLER_0_12_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08053_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09368__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08142__C team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1119_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout481_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _03789_ _03792_ _03772_ _03781_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08886_ net1551 _04573_ _04557_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
X_16722__1276 vssd1 vssd1 vccd1 vccd1 _16722__1276/HI net1276 sky130_fd_sc_hd__conb_1
XANTENNA__09540__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _03685_ _03724_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07768_ _03611_ _03651_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\] net812 net848 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15575__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _03586_ _03589_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout913_A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11305__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09438_ net609 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[21\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09369_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] net652 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11400_ net454 _06146_ _07007_ net438 _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12060__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12380_ net306 net1870 net495 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ net417 _06508_ _06944_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14050_ net1090 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XANTENNA__09359__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11262_ net450 _06877_ _06879_ _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13001_ net229 _03024_ _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__nand3_1
X_10213_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] net651 _05868_ vssd1
+ vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a21o_1
XANTENNA__12570__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ net393 _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__and2_1
XANTENNA_input42_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\] net842 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14952_ net1195 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
X_10075_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] net766 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\]
+ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__a221o_1
XANTENNA__10126__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ net1125 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
X_14883_ net1158 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XANTENNA__15918__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11914__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16622_ clknet_leaf_65_wb_clk_i _02856_ _01495_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_13834_ net1050 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13765_ net1075 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
X_16553_ clknet_leaf_5_wb_clk_i net1418 _01426_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10977_ _06611_ _06612_ net909 vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and3b_1
X_15504_ clknet_leaf_34_wb_clk_i _01955_ _00462_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12716_ team_02_WB.instance_to_wrap.top.i_ready _04513_ _07335_ team_02_WB.instance_to_wrap.top.pc\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16484_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[19\] _01358_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[19\] sky130_fd_sc_hd__dfrtp_1
X_13696_ net1078 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15435_ clknet_leaf_21_wb_clk_i _01886_ _00393_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12647_ _04743_ _04784_ _06135_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ clknet_leaf_12_wb_clk_i _01817_ _00324_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12578_ net303 net2304 net475 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14317_ net1134 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
X_11529_ _06006_ _06159_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__xor2_1
X_15297_ clknet_leaf_130_wb_clk_i _01748_ _00255_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold307 team_02_WB.instance_to_wrap.top.pc\[3\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold318 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold329 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1083 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12480__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ net1069 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout809 _04657_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__buf_6
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09770__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11096__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1007 net113 vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_08740_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[22\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[22\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_2
Xhold1018 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08671_ net745 _04449_ _04455_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__and3_4
XANTENNA__15598__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11824__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03510_ _03511_ _03512_ vssd1
+ vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07553_ _03435_ _03437_ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1
+ vccd1 vccd1 _03444_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07484_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] net1689 net964 vssd1
+ vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\] net816 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1069_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09589__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ _04828_ _04830_ _04832_ _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__or4_2
XFILLER_0_8_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08105_ _03971_ _03975_ _03982_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__o31a_1
XANTENNA__08797__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] net870 net794 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\]
+ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08036_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
Xhold830 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold841 team_02_WB.instance_to_wrap.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net2239
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12390__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07484__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09761__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\] net791 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout863_A _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08938_ _04616_ _04618_ _04620_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__or4_2
XFILLER_0_99_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11856__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08869_ net1557 _04562_ net825 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__mux2_1
X_10900_ _06209_ _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__or2_1
XANTENNA__11734__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880_ net295 net2223 net544 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08609__A team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _06475_ _06477_ _06478_ team_02_WB.instance_to_wrap.top.aluOut\[29\] net460
+ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__o32a_4
XFILLER_0_95_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13234__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16826__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _03387_ _03388_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10762_ _04625_ net401 vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ net2427 net243 net478 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10831__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] _03342_ vssd1 vssd1 vccd1
+ vccd1 _03343_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10874__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ team_02_WB.instance_to_wrap.top.pc\[30\] team_02_WB.instance_to_wrap.top.pc\[29\]
+ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15220_ clknet_leaf_53_wb_clk_i _01671_ _00178_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ net233 net1764 net490 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__mux2_1
XANTENNA__10593__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15151_ clknet_leaf_32_wb_clk_i _01602_ _00109_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12363_ net354 net2186 net499 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14102_ net1105 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ team_02_WB.instance_to_wrap.top.pc\[12\] _06333_ team_02_WB.instance_to_wrap.top.pc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15082_ clknet_leaf_77_wb_clk_i _01533_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.halfData\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12294_ net337 net2700 net505 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11909__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14033_ net1028 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ _05379_ _05397_ _06865_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10898__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _05235_ net431 net447 _05237_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10127_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] net799 _05783_ _05785_
+ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__a211o_1
X_15984_ clknet_leaf_39_wb_clk_i _02435_ _00942_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09504__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10058_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] net709 net702 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a221o_1
X_14935_ net1008 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11644__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14866_ net1171 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ clknet_leaf_61_wb_clk_i _02839_ _01478_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_13817_ net1064 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14797_ net1198 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_69_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16536_ clknet_leaf_0_wb_clk_i net1446 _01409_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ net1038 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10822__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16467_ clknet_leaf_99_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[2\] _01341_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[2\] sky130_fd_sc_hd__dfrtp_1
X_13679_ net1127 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XANTENNA__14256__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12024__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15418_ clknet_leaf_120_wb_clk_i _01869_ _00376_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11599__B _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16398_ clknet_leaf_78_wb_clk_i net1464 _01272_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.flip2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08779__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16721__1275 vssd1 vssd1 vccd1 vccd1 _16721__1275/HI net1275 sky130_fd_sc_hd__conb_1
XFILLER_0_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ clknet_leaf_116_wb_clk_i _01800_ _00307_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 _02586_ vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10050__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold115 _02598_ vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09991__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1
+ net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1 net1535
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _02590_ vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11819__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] net661 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a22o_1
Xhold159 team_02_WB.instance_to_wrap.top.a1.data\[7\] vssd1 vssd1 vccd1 vccd1 net1557
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10338__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] net856 net756 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\]
+ _05504_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a221o_1
Xfanout617 net619 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09743__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout628 net631 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_8
Xfanout639 _04488_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09772_ _05432_ _05434_ _05436_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__or4_1
XANTENNA__13288__C1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08723_ net1654 net955 net926 _04518_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16631__1379 vssd1 vssd1 vccd1 vccd1 net1379 _16631__1379/LO sky130_fd_sc_hd__conb_1
X_08654_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] net731 net726 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _03453_ _03465_ _03472_ _03457_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08585_ _04379_ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout444_A _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1186_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] _03426_ vssd1 vssd1 vccd1
+ vccd1 _03427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08863__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12893__B _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07467_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 _03407_
+ sky130_fd_sc_hd__inv_2
XANTENNA__12385__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout709_A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07479__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\] net645 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\]
+ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15613__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] net858 net850 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] net674 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a22o_1
XANTENNA__09982__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08019_ _03902_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nand2_1
XANTENNA__11729__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15763__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold671 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net441 _06647_ _06666_ net428 _06662_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[23\]
+ sky130_fd_sc_hd__a221o_2
Xhold693 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07508__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12981_ _06614_ _07335_ _02966_ _03004_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13245__A team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14720_ net1040 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ net358 net2303 net540 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14651_ net1043 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
X_11863_ net342 net2211 net548 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XANTENNA__13046__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13602_ net1087 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
X_10814_ net400 _06462_ _06424_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__o21a_1
XANTENNA__11057__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11057__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14582_ net1111 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
X_11794_ net337 net2733 net557 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16321_ clknet_leaf_96_wb_clk_i _02754_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13533_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] _03376_
+ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__and2_1
X_10745_ _06388_ _06395_ net390 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12295__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15293__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13464_ net1641 _03331_ _03333_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__o21a_1
X_16252_ clknet_leaf_98_wb_clk_i _02690_ _01209_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10676_ team_02_WB.instance_to_wrap.top.pc\[4\] team_02_WB.instance_to_wrap.top.pc\[3\]
+ team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12415_ net321 net1807 net490 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15203_ clknet_leaf_42_wb_clk_i _01654_ _00161_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16183_ clknet_leaf_66_wb_clk_i _02629_ _01141_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13395_ team_02_WB.instance_to_wrap.top.a1.row2\[15\] _03206_ _03280_ _03273_ team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10032__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12346_ net295 net2445 net496 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__mux2_1
X_15134_ clknet_leaf_5_wb_clk_i _01585_ _00092_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11639__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15065_ clknet_leaf_59_wb_clk_i _01516_ _00028_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[18\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_116_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12277_ net273 net1882 net505 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14016_ net1078 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
X_11228_ net419 _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__nor2_1
XANTENNA__09725__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ _05238_ _06030_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15967_ clknet_leaf_9_wb_clk_i _02418_ _00925_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14918_ net1164 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15898_ clknet_leaf_120_wb_clk_i _02349_ _00856_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14849_ net1155 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08370_ _04243_ _04239_ _04236_ _04235_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__15636__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09110__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16519_ clknet_leaf_5_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[22\]
+ _01393_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10271__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15786__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10023__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09177__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout403 net406 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
XANTENNA__09716__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_2
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 _06120_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08924__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09824_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\] net683 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a22o_1
Xfanout447 _06134_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_2
Xfanout458 _06326_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1101_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net471 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_4
XANTENNA__12888__B _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15166__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\] net865 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__a22o_1
XANTENNA__10689__A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16411__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04367_ _04426_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a22o_1
XANTENNA__11287__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11287__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ _05349_ _05352_ _05353_ _05354_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[15\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_90_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08637_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13028__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08568_ net973 net975 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16561__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ net1825 _03414_ net1 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16526__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08499_ team_02_WB.instance_to_wrap.top.a1.row1\[61\] _04333_ _04325_ vssd1 vssd1
+ vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10530_ _06154_ _06169_ _06170_ _06182_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10262__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12200_ net234 net2313 net519 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13180_ _03144_ _03163_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o21a_1
XANTENNA__09955__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ _06042_ _06044_ _04952_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__o21a_1
X_12131_ net357 net2696 net589 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
XANTENNA__11459__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ net340 net2422 net530 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09707__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15509__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11013_ _06534_ _06649_ net384 vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08768__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_2
XFILLER_0_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_1
X_15821_ clknet_leaf_23_wb_clk_i _02272_ _00779_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16720__1274 vssd1 vssd1 vccd1 vccd1 _16720__1274/HI net1274 sky130_fd_sc_hd__conb_1
X_15752_ clknet_leaf_56_wb_clk_i _02203_ _00710_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12964_ _02883_ _02969_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1190 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09340__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14703_ net1169 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
X_11915_ net316 net1967 net542 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ clknet_leaf_45_wb_clk_i _02134_ _00641_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ team_02_WB.instance_to_wrap.top.pc\[2\] _05936_ vssd1 vssd1 vccd1 vccd1 _02929_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__08694__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13703__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ net1162 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ net287 net2131 net548 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14565_ net1076 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11777_ net271 net1881 net559 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XANTENNA__10789__B1 team_02_WB.instance_to_wrap.top.aluOut\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16304_ clknet_leaf_80_wb_clk_i _02737_ _01247_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13516_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1
+ vccd1 _03366_ sky130_fd_sc_hd__and3_1
X_10728_ _06375_ _06378_ net363 vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__mux2_1
XANTENNA__10253__A2 _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14496_ net1071 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16235_ clknet_leaf_78_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] _01192_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[3\] sky130_fd_sc_hd__dfrtp_1
X_10659_ team_02_WB.instance_to_wrap.top.pc\[28\] _06229_ _06310_ vssd1 vssd1 vccd1
+ vccd1 _06311_ sky130_fd_sc_hd__a21o_1
X_13447_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] _03321_ net1175 vssd1 vssd1
+ vccd1 vccd1 _03323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14534__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10005__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ clknet_leaf_71_wb_clk_i _02612_ _01124_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09946__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630__1378 vssd1 vssd1 vccd1 vccd1 net1378 _16630__1378/LO sky130_fd_sc_hd__conb_1
X_13378_ team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] _03217_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15117_ clknet_leaf_24_wb_clk_i _01568_ _00075_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12329_ net344 net2175 net502 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16097_ clknet_leaf_92_wb_clk_i _02543_ _01055_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09159__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15048_ net1164 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__inv_2
XANTENNA__15189__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07870_ _03729_ _03757_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\] net677 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09471_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] net805 net793 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\]
+ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a221o_1
XANTENNA__09882__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08685__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09882__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14709__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11832__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12218__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08422_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[11\] _04277_ vssd1 vssd1 vccd1
+ vccd1 _04287_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07611__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ net1719 net935 net918 _04228_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10448__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08437__A2 _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10244__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__A1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08284_ _04140_ _04151_ _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_127_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11279__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout776_A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout233 net236 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net257 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09570__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _06618_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
X_09807_ _05469_ _05470_ _05471_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__or4_1
Xfanout288 net290 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlymetal6s2s_1
X_07999_ _03856_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 net302 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net728 net676 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09322__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09669_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\] net805 net797 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11742__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15951__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ net234 net1747 net569 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ _06744_ _06877_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__or2_1
XANTENNA__10483__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ net358 net1846 net576 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XANTENNA__13242__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14350_ net1063 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XANTENNA__10235__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ net366 _06108_ _06111_ net386 vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08055__C _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ _05722_ _05746_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__o21ai_1
X_13301_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] _03206_ vssd1 vssd1 vccd1
+ vccd1 _03207_ sky130_fd_sc_hd__nand2_1
X_14281_ net1007 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XANTENNA__12573__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] net887 net907 team_02_WB.instance_to_wrap.top.pc\[5\]
+ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16020_ clknet_leaf_47_wb_clk_i _02471_ _00978_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13232_ team_02_WB.instance_to_wrap.ramload\[5\] net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[5\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09389__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _05591_ net368 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__nand2_1
XANTENNA_input72_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15331__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13163_ team_02_WB.instance_to_wrap.top.lcd.currentState\[1\] net986 net895 vssd1
+ vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10375_ _05257_ _05275_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10943__B1 _06569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12114_ net297 net2526 net586 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13094_ team_02_WB.instance_to_wrap.top.pc\[7\] net946 net941 _03103_ vssd1 vssd1
+ vccd1 vccd1 _01505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11917__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ net271 net1772 net530 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09561__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15804_ clknet_leaf_49_wb_clk_i _02255_ _00762_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16784_ net1338 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996_ net1003 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ clknet_leaf_119_wb_clk_i _02186_ _00693_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12947_ _02973_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11120__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08667__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11652__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15666_ clknet_leaf_10_wb_clk_i _02117_ _00624_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12878_ _02911_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14617_ net1164 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ net344 net2076 net554 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__mux2_1
X_15597_ clknet_leaf_43_wb_clk_i _02048_ _00555_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11423__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ net1052 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09092__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12483__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14479_ net1124 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16218_ clknet_leaf_35_wb_clk_i _02663_ _01175_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09919__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ clknet_leaf_129_wb_clk_i net1531 _01107_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15824__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ net972 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ net886 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__o31a_2
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11827__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _03810_ _03811_ _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a21bo_1
Xhold19 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[30\] vssd1 vssd1 vccd1 vccd1
+ net1417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09552__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _03703_ _03737_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07606__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15974__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _03642_ _03673_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09304__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout357_A _07135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\] net736 net688 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1099_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15204__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10686__B team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08405_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ team_02_WB.instance_to_wrap.top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_34_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] net855 net781 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout524_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10217__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08336_ _04189_ _04191_ _04196_ _04190_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08871__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15354__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ _04121_ _04136_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08830__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08198_ _04073_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10160_ net897 _05797_ _05815_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09791__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11737__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1015 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1017 net1019 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
X_10091_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\] net709 net661 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__a22o_1
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_4
Xfanout1039 net1049 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13850_ net1052 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08897__A_N net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12801_ _07407_ _07422_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__o21a_1
XANTENNA__09731__A _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13781_ net1114 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XANTENNA__12568__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _06563_ _06631_ net379 vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__mux2_1
XANTENNA__14349__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15520_ clknet_leaf_9_wb_clk_i _01971_ _00478_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12732_ _07353_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15451_ clknet_leaf_104_wb_clk_i _01902_ _00409_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12663_ _07272_ _07282_ _07283_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14402_ net1088 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
X_11614_ net316 net2540 net578 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XANTENNA__10208__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15382_ clknet_leaf_108_wb_clk_i _01833_ _00340_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09074__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ net355 net2190 net475 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ net1031 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
X_11545_ _05863_ _06981_ _07139_ net411 vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__o211a_1
XANTENNA__14084__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14264_ net1114 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
X_11476_ _05837_ _06008_ _06011_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__nor3_1
XANTENNA__15847__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16003_ clknet_leaf_45_wb_clk_i _02454_ _00961_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13215_ team_02_WB.START_ADDR_VAL_REG\[23\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net207 sky130_fd_sc_hd__a21o_1
X_10427_ _06078_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14195_ net1127 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XANTENNA__14812__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13146_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__and4bb_1
X_10358_ _05793_ _06009_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16815__1369 vssd1 vssd1 vccd1 vccd1 _16815__1369/HI net1369 sky130_fd_sc_hd__conb_1
XFILLER_0_57_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11647__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15997__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ team_02_WB.instance_to_wrap.top.pc\[10\] net945 net941 _03089_ vssd1 vssd1
+ vccd1 vccd1 _01508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10289_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\] net821 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ _05937_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09534__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ net336 net1761 net468 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
XANTENNA__07545__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12478__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ net1321 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
XANTENNA__13094__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13979_ net1045 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XANTENNA__10787__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15718_ clknet_leaf_11_wb_clk_i _02169_ _00676_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16698_ net1252 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15377__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15649_ clknet_leaf_1_wb_clk_i _02100_ _00607_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\] net806 net778 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09065__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ _03993_ _03996_ _03998_ _04000_ _03992_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__o311a_1
XFILLER_0_56_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08052_ _03937_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08954_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ net886 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__and3b_2
XANTENNA_fanout1014_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _03780_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__nor2_1
X_08885_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] net939 _04571_ _04572_ vssd1
+ vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout474_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07836_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] _03724_ _03725_ vssd1 vssd1
+ vccd1 vccd1 _03727_ sky130_fd_sc_hd__or3_1
XANTENNA__12896__B _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12388__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _03611_ _03651_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout641_A _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout739_A _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[19\] net859 net767 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\]
+ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07698_ _03587_ _03588_ _03544_ net362 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09437_ _05098_ _05107_ _05110_ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__nor4_1
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] net726 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__a221o_1
XANTENNA__09056__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11399__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ _04194_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__nand2_1
X_09299_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] net767 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08803__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10071__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ net417 _06507_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__a21o_1
XANTENNA__10522__A_N _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11261_ _05359_ net433 _06880_ _06056_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10212_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\] net739 net683 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a22o_1
X_13000_ _02892_ _02893_ _02961_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__nand3_1
XANTENNA__09764__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _06709_ _06816_ net382 vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10143_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\] net785 net781 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\]
+ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a221o_1
XANTENNA__09516__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A wbm_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ net1047 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
X_10074_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] net871 net862 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13902_ net1116 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
X_14882_ net1150 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XANTENNA__08776__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ clknet_leaf_60_wb_clk_i _02855_ _01494_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09461__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ net1012 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XANTENNA__12298__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16552_ clknet_leaf_5_wb_clk_i net1413 _01425_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13764_ net1142 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
X_10976_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net744 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ net443 vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__a221o_1
XANTENNA__09295__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15503_ clknet_leaf_32_wb_clk_i _01954_ _00461_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ net231 _07331_ _07332_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16483_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[18\] _01357_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13695_ net1130 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11930__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15434_ clknet_leaf_46_wb_clk_i _01885_ _00392_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12646_ _04825_ _04867_ _04912_ _04952_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__or4_1
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09047__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15365_ clknet_leaf_127_wb_clk_i _01816_ _00323_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08255__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ net295 net1822 net472 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
X_14316_ net1006 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ net419 _06766_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ clknet_leaf_6_wb_clk_i _01747_ _00254_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold308 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ net1136 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
X_11459_ _06980_ _07061_ net386 vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09755__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ net1090 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XANTENNA__11562__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ _00006_ team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] vssd1 vssd1 vccd1
+ vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] sky130_fd_sc_hd__or2_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09507__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1019 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ net745 _04454_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__and3_4
XFILLER_0_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07533__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ _03476_ _03506_ _03406_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16819_ net1373 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XFILLER_0_17_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07552_ _03428_ _03435_ _03442_ _03405_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12001__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09286__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07483_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] team_02_WB.instance_to_wrap.ramload\[22\]
+ net964 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14717__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11840__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[26\] net796 net790 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\]
+ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08715__A _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09153_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] net684 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08104_ _03984_ _03986_ _03989_ _03983_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__o22a_1
XANTENNA__10053__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] net843 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08035_ _03863_ _03895_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput80 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold820 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput91 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold831 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold842 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09746__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16518__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold864 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold886 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A _04468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold897 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\] net815 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08937_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[31\] net732 net696 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[31\]
+ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout856_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15542__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ net959 _04300_ _04311_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07819_ _03686_ _03687_ _03682_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a21o_2
X_08799_ net166 net951 net903 net1496 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08609__B team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10830_ _06225_ net744 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[29\] net443
+ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15692__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ _04625_ net421 vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__nand2_2
XANTENNA__08485__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11750__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ net2622 net239 net478 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16814__1368 vssd1 vssd1 vccd1 vccd1 _16814__1368/HI net1368 sky130_fd_sc_hd__conb_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ team_02_WB.instance_to_wrap.top.pc\[28\] team_02_WB.instance_to_wrap.top.pc\[27\]
+ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__and3_1
XANTENNA__09029__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13480_ net873 _03341_ _03342_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16048__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08237__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ net358 net1949 net488 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__mux2_1
XANTENNA__10044__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ clknet_leaf_40_wb_clk_i _01601_ _00108_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09985__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net344 net2101 net496 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14101_ net1118 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11313_ _06274_ _06277_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__nand2_1
X_15081_ clknet_leaf_78_wb_clk_i _01532_ _00044_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_12293_ net334 net2538 net504 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XANTENNA__12581__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14032_ net1016 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XANTENNA__09737__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ _05402_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09201__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11175_ net435 _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__nor2_1
X_10126_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net811 net787 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a221o_1
X_15983_ clknet_leaf_33_wb_clk_i _02434_ _00941_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11925__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] net718 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a22o_1
X_14934_ net1034 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XANTENNA__08712__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08712__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ net1171 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16604_ clknet_leaf_61_wb_clk_i _02838_ _01477_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13816_ net1107 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
XANTENNA__09268__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14796_ net1198 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16535_ clknet_leaf_1_wb_clk_i net1426 _01408_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08476__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ net1128 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
X_10959_ net384 _06599_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11660__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10283__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16466_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[1\] _01340_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13678_ net1116 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15417_ clknet_leaf_108_wb_clk_i _01868_ _00375_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ _07252_ _07253_ _07254_ _07256_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__or4b_1
X_16397_ clknet_leaf_78_wb_clk_i team_02_WB.instance_to_wrap.top.edg2.button_i _01271_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.flip1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10035__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08779__B2 _04546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15415__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15348_ clknet_leaf_51_wb_clk_i _01799_ _00306_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12491__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[20\] vssd1 vssd1 vccd1
+ vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15279_ clknet_leaf_31_wb_clk_i _01730_ _00237_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold116 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[2\] vssd1 vssd1 vccd1
+ vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 team_02_WB.instance_to_wrap.top.a1.row1\[108\] vssd1 vssd1 vccd1 vccd1 net1525
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[14\] vssd1 vssd1 vccd1
+ vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net1547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11535__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09840_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\] net881 net877 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08400__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_8
Xfanout629 net631 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_4
XFILLER_0_123_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] net809 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08722_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[31\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[31\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09900__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ net747 _04443_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__and3_4
XANTENNA__10510__A1 _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ _03464_ _03491_ _03492_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09259__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ _03396_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07535_ team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] team_02_WB.instance_to_wrap.top.a1.dataIn\[20\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1 vccd1 _03426_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10975__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 _03406_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_107_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08445__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08482__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] net662 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a22o_1
XANTENNA__10026__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] net767 net838 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a221o_1
XANTENNA__09967__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] net713 _04749_ vssd1
+ vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15908__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07495__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09719__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03903_ _03904_ _03905_ vssd1
+ vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold650 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold672 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold694 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14910__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09969_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\] net709 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a221o_1
XANTENNA__11745__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ _03006_ _03007_ _04514_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09498__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1350 team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net2748
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11931_ net351 net2147 net540 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14650_ net1003 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
X_11862_ net349 net2257 net549 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ net1102 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10813_ net388 _06461_ _06421_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14581_ net1117 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XANTENNA__12576__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net335 net2521 net556 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10265__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16320_ clknet_leaf_97_wb_clk_i _02753_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13532_ _03376_ net885 _03375_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__and3b_1
XFILLER_0_113_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15438__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10744_ _06391_ _06394_ net366 vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09670__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16251_ clknet_leaf_93_wb_clk_i _02689_ _01208_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_13463_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] _03331_ net1176 vssd1
+ vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__a21oi_1
X_10675_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net744 net458 team_02_WB.instance_to_wrap.top.a1.dataIn\[31\]
+ net444 vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15202_ clknet_leaf_49_wb_clk_i _01653_ _00160_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12414_ net317 net2589 net489 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16182_ clknet_leaf_71_wb_clk_i _02628_ _01140_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13394_ _03206_ _03281_ _03291_ _03292_ _03142_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09422__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15588__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ clknet_leaf_117_wb_clk_i _01584_ _00091_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ net287 net1753 net496 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15064_ clknet_leaf_59_wb_clk_i _01515_ _00027_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_12276_ net277 net2144 net506 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11517__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12714__C1 team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09186__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ net1131 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
X_11227_ _06633_ _06849_ net397 vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__mux2_1
XANTENNA__14820__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11158_ _06293_ _06784_ net909 vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and3b_1
XANTENNA__11655__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10109_ _05758_ _05767_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nor2_4
X_15966_ clknet_leaf_12_wb_clk_i _02417_ _00924_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11089_ team_02_WB.instance_to_wrap.top.pc\[21\] _06339_ vssd1 vssd1 vccd1 vccd1
+ _06721_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09489__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10390__A_N _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ net1165 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XANTENNA__08697__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ clknet_leaf_117_wb_clk_i _02348_ _00855_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14848_ net1155 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12994__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12486__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14779_ net1177 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16652__1219 vssd1 vssd1 vccd1 vccd1 _16652__1219/HI net1219 sky130_fd_sc_hd__conb_1
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10256__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16518_ clknet_leaf_5_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[21\]
+ _01392_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16363__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08265__A team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09661__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16449_ clknet_leaf_82_wb_clk_i net1469 _01323_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09413__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07975__A2 _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 net406 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
Xfanout415 _05817_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
X_09823_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] net687 net643 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[11\]
+ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a221o_1
X_16813__1367 vssd1 vssd1 vccd1 vccd1 _16813__1367/HI net1367 sky130_fd_sc_hd__conb_1
Xfanout437 _06057_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 _06132_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 _04582_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _05411_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nor2_8
XFILLER_0_20_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08705_ _04473_ _04498_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nor2_4
XANTENNA__08688__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] net878 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ _05339_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08636_ _04402_ _04430_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07998__B _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net973 net975 vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10247__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07518_ net2390 net991 net2 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08498_ net940 _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__or2_1
XANTENNA__09652__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ _06111_ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09404__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net717 net674 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10391_ _04991_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12130_ net345 net1981 net588 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
XANTENNA__15880__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ net336 net2516 net528 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold480 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold491 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012_ _06598_ _06648_ net378 vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__mux2_1
XANTENNA__09734__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12784__A_N _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15820_ clknet_leaf_52_wb_clk_i _02271_ _00778_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout960 _04272_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_2
Xfanout971 _03413_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 net984 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15751_ clknet_leaf_15_wb_clk_i _02202_ _00709_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12963_ _02993_ _02991_ _07364_ team_02_WB.instance_to_wrap.top.pc\[28\] vssd1 vssd1
+ vccd1 vccd1 _01526_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08679__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1180 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ net1167 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
Xhold1191 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ net303 net1973 net543 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
X_15682_ clknet_leaf_47_wb_clk_i _02133_ _00640_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15260__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08784__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ team_02_WB.instance_to_wrap.top.pc\[3\] _05889_ vssd1 vssd1 vccd1 vccd1 _02928_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ net1158 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
X_11845_ net282 net1837 net549 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14087__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10238__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14564_ net1145 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
X_11776_ net277 net1792 net558 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09643__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10789__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16303_ clknet_leaf_92_wb_clk_i _02736_ _01246_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13515_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] net1690
+ _03365_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a21oi_1
X_10727_ _06376_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__nand2_1
XANTENNA__08851__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14495_ net1121 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XANTENNA__11450__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14815__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16234_ clknet_leaf_78_wb_clk_i _00006_ _01191_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13446_ _03321_ _03322_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__nor2_1
X_10658_ _06230_ _06309_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16165_ clknet_leaf_66_wb_clk_i _02611_ _01123_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13377_ team_02_WB.instance_to_wrap.top.a1.row1\[12\] _03217_ _03221_ _03226_ team_02_WB.instance_to_wrap.top.a1.row1\[60\]
+ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a32o_1
X_10589_ team_02_WB.instance_to_wrap.top.a1.instruction\[24\] net928 net590 vssd1
+ vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__a21oi_4
X_15116_ clknet_leaf_52_wb_clk_i _01567_ _00074_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ net348 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\] net502 vssd1
+ vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
X_16096_ clknet_leaf_92_wb_clk_i _02542_ _01054_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ net1164 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__inv_2
X_12259_ net330 net1721 net510 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12989__B _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15603__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15949_ clknet_leaf_24_wb_clk_i _02400_ _00907_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09470_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\] net821 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08005__A2_N _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ team_02_WB.instance_to_wrap.top.a1.state\[1\] _04284_ _04286_ net1736 vssd1
+ vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ _04220_ _04225_ _04227_ _04217_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09634__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08842__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ _04145_ _04149_ _04150_ _04142_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13194__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout302_A _06956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08869__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout671_A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout245 _06439_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout769_A _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\] net779 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\]
+ _05463_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a221o_1
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
Xfanout278 _06645_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15283__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ _03851_ _03860_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__nand2_2
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] net716 net704 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09668_ _05327_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__nor2_8
XFILLER_0_35_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09873__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08619_ net977 net931 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nand2b_4
X_09599_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\] net767 _05259_ _05261_
+ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11630_ net352 net2045 net576 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XANTENNA__09086__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__B1 _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08833__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11561_ net365 _07120_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__nand2_1
Xwire602 _05654_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire613 _04822_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
X_13300_ _03398_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] vssd1 vssd1 vccd1
+ vccd1 _03206_ sky130_fd_sc_hd__nor2_2
X_10512_ _05749_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14280_ net1083 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11492_ net913 _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ team_02_WB.instance_to_wrap.ramload\[4\] net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[4\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ _06094_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input65_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13162_ net992 _03151_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10374_ _05318_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10943__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ net290 net2386 net586 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XANTENNA__14370__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _07428_ _03101_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__o21ai_1
X_16651__1218 vssd1 vssd1 vccd1 vccd1 _16651__1218/HI net1218 sky130_fd_sc_hd__conb_1
X_12044_ net276 net2492 net529 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net792 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15803_ clknet_leaf_119_wb_clk_i _02254_ _00761_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16783_ net1337 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
X_13995_ net1030 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11933__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15734_ clknet_leaf_111_wb_clk_i _02185_ _00692_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12946_ _02876_ _02877_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09864__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11120__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15665_ clknet_leaf_111_wb_clk_i _02116_ _00623_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12877_ team_02_WB.instance_to_wrap.top.pc\[12\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _02911_ sky130_fd_sc_hd__and2_1
X_14616_ net1156 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09077__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ net347 net2359 net554 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__mux2_1
X_15596_ clknet_leaf_52_wb_clk_i _02047_ _00554_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547_ net1128 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
X_16812__1366 vssd1 vssd1 vccd1 vccd1 _16812__1366/HI net1366 sky130_fd_sc_hd__conb_1
X_11759_ net330 net2683 net561 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478_ net1117 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15156__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16217_ clknet_leaf_38_wb_clk_i _02662_ _01174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13429_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _03312_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16148_ clknet_leaf_6_wb_clk_i net1569 _01106_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16079_ clknet_leaf_35_wb_clk_i _02530_ _01037_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_08970_ net883 _04637_ _04651_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_100_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12136__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07921_ _03765_ _03766_ _03789_ _03792_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09001__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12004__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _03742_ _03741_ _03693_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__and3b_1
XANTENNA__07563__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_07783_ _03642_ _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11843__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09522_ _05175_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09453_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[20\] net712 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout252_A _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ net990 net991 _04269_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] vssd1
+ vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__or4b_1
XFILLER_0_8_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09068__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] net797 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ _04199_ _04200_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08815__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout517_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08266_ _04121_ _04136_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nand2_1
XANTENNA__08453__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08197_ _04048_ _04076_ _04077_ _04078_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or4_1
XANTENNA__11178__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11178__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15649__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout886_A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ _05747_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__nor2_2
Xfanout1007 net1010 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_4
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_4
Xfanout1029 net1032 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15799__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11753__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _07406_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__nor2_1
X_13780_ net1036 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_10992_ _06373_ _06377_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__nand2_1
XANTENNA__09846__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08628__A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ _03418_ _03420_ _07357_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15450_ clknet_leaf_120_wb_clk_i _01901_ _00408_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12662_ _05701_ _05747_ _07288_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ net1102 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
X_11613_ net303 net2374 net578 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15381_ clknet_leaf_115_wb_clk_i _01832_ _00339_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12584__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08806__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16424__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ net342 net1970 net473 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__mux2_1
XANTENNA__10893__A _06132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ net1102 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_11544_ net392 _07061_ _07138_ net404 vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ net1115 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
X_11475_ _06011_ _06162_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16002_ clknet_leaf_47_wb_clk_i _02453_ _00960_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13214_ team_02_WB.START_ADDR_VAL_REG\[22\] _04356_ vssd1 vssd1 vccd1 vccd1 net206
+ sky130_fd_sc_hd__and2_1
XFILLER_0_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10426_ _04888_ net373 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14194_ net1085 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11928__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _03138_
+ sky130_fd_sc_hd__or3b_1
XANTENNA__10832__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10357_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__inv_2
XANTENNA__12118__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13076_ net230 _03086_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__a21bo_1
X_10288_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] net801 net785 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\]
+ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12027_ net333 net2125 net469 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
XANTENNA__10144__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__B2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11663__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13978_ net1045 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09298__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ net1320 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XFILLER_0_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15717_ clknet_leaf_125_wb_clk_i _02168_ _00675_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12929_ _02892_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16697_ net1251 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ clknet_leaf_6_wb_clk_i _02099_ _00606_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13397__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15579_ clknet_leaf_106_wb_clk_i _02030_ _00537_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ _03971_ _03975_ _03982_ _04002_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o31a_2
XFILLER_0_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08051_ _03902_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09222__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08953_ net883 _04636_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07876__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ _03790_ _03791_ _03771_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08884_ net959 _04318_ _04328_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1
+ vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a22o_1
X_07835_ _03724_ _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout467_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07766_ _03655_ _03656_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nor2_2
XANTENNA__09289__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09505_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] net852 net832 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07697_ _03510_ _03542_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__A team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] net849 net777 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[21\]
+ _05096_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08882__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13388__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16650__1217 vssd1 vssd1 vccd1 vccd1 _16650__1217/HI net1217 sky130_fd_sc_hd__conb_1
X_09367_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\] net738 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout801_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07498__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08318_ _04181_ _04182_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__nand2_2
XFILLER_0_62_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09298_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[24\] net846 net838 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08249_ _04103_ _04119_ _04104_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11260_ _05357_ net446 _06151_ net455 vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09213__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13014__A1_N net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] net735 net707 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a221o_1
XANTENNA__11748__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11191_ _06760_ _06815_ net376 vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11571__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10142_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] net817 net761 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a22o_1
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 wbm_we_o sky130_fd_sc_hd__buf_2
XFILLER_0_105_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14950_ net1034 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
X_10073_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] net795 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a221o_1
XANTENNA__10126__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16811__1365 vssd1 vssd1 vccd1 vccd1 _16811__1365/HI net1365 sky130_fd_sc_hd__conb_1
X_13901_ net1132 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XANTENNA_input28_A wbm_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1150 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XANTENNA__12579__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16620_ clknet_leaf_62_wb_clk_i _02854_ _01493_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_13832_ net1096 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XANTENNA__13076__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16551_ clknet_leaf_129_wb_clk_i net1448 _01424_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13763_ net1068 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ net911 _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15502_ clknet_leaf_42_wb_clk_i _01953_ _00460_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12714_ net889 _07340_ _07341_ net228 team_02_WB.instance_to_wrap.top.i_ready vssd1
+ vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__o311ai_1
X_16482_ clknet_leaf_75_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[17\] _01356_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[17\] sky130_fd_sc_hd__dfrtp_1
X_13694_ net1020 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15814__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15433_ clknet_leaf_29_wb_clk_i _01884_ _00391_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12645_ _05702_ _05748_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15364_ clknet_leaf_53_wb_clk_i _01815_ _00322_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09189__A _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ net288 net1763 net472 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14315_ net1014 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
X_11527_ net394 _06961_ _07122_ _07123_ net408 vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15964__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15295_ clknet_leaf_26_wb_clk_i _01746_ _00253_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold309 team_02_WB.instance_to_wrap.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net1707
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ net1092 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09204__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ _07020_ _07060_ net381 vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11658__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _05296_ net372 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14177_ net1143 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ _05656_ _06015_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__and2b_1
X_13128_ _04270_ net1677 _03126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[1\]
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13059_ _06954_ net227 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__or2_1
Xhold1009 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15344__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12489__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07620_ _03406_ _03506_ _03476_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a21boi_1
XANTENNA__13174__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16818_ net1372 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07551_ _03435_ _03437_ _03426_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16749_ net1303 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07482_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] net2728 net964 vssd1
+ vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\] net802 net770 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\] net733 net721 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09443__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08103_ _03983_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__or2_2
XANTENNA__09994__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] net818 net754 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14733__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08034_ _03912_ _03921_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput70 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_1
Xhold810 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput81 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold821 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput92 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
Xhold832 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 team_02_WB.instance_to_wrap.ramload\[7\] vssd1 vssd1 vccd1 vccd1 net2241
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16370__D _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold854 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold865 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold898 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09985_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] net867 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout584_A _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net716 net700 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08867_ net1575 _04561_ net825 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__mux2_1
XANTENNA__12399__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout849_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _03698_ _03706_ _03707_ _03703_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__or4b_2
X_08798_ net167 net952 net903 net1471 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XANTENNA__13058__B2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15837__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ _03577_ _03638_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14908__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10760_ net580 net414 vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__nor2_1
XANTENNA__09682__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09419_ _05084_ _05093_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nor2_4
X_10691_ team_02_WB.instance_to_wrap.top.pc\[26\] _06342_ vssd1 vssd1 vccd1 vccd1
+ _06343_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15987__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12430_ net353 net2038 net488 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09434__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ net348 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\] net498 vssd1
+ vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14100_ net1051 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
X_11312_ net426 _06914_ _06928_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[13\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15080_ clknet_leaf_78_wb_clk_i _01531_ _00043_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12292_ net330 net2108 net505 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08641__A team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14031_ net1125 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11243_ _06176_ _06863_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ net417 _06794_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__or2_1
XANTENNA__15367__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] net859 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__a22o_1
XANTENNA__16612__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ clknet_leaf_40_wb_clk_i _02433_ _00940_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10056_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] net738 net698 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\]
+ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a221o_1
X_14933_ net1010 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11507__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14864_ net1172 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
X_16603_ clknet_leaf_60_wb_clk_i _02837_ _01476_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13815_ net1107 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14795_ net1174 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11941__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16534_ clknet_leaf_36_wb_clk_i net1414 _01407_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13746_ net1082 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
X_10958_ _06533_ _06598_ net378 vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__mux2_1
XANTENNA__09673__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ net1135 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16465_ clknet_leaf_81_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[0\] _01339_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[0\] sky130_fd_sc_hd__dfrtp_1
X_10889_ _06460_ _06533_ net378 vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15416_ clknet_leaf_121_wb_clk_i _01867_ _00374_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12628_ _06759_ _06846_ _07255_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__and3_1
X_16396_ clknet_leaf_74_wb_clk_i _02827_ _01270_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09425__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ clknet_leaf_124_wb_clk_i _01798_ _00305_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11232__B1 _06846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ net346 net2082 net465 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12980__B1 _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__A _05296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ clknet_leaf_39_wb_clk_i _01729_ _00236_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold106 _02599_ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 _02581_ vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold128 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[28\] vssd1 vssd1 vccd1
+ vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14229_ net1115 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
Xhold139 _02593_ vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11535__A1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10338__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08400__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout619 _04496_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09770_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\] net869 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13288__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08721_ net988 _03404_ _04341_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_4
X_08652_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and3b_2
XANTENNA__12012__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ _03453_ _03465_ _03472_ _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__o31ai_2
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04367_ vssd1 vssd1 vccd1
+ vccd1 _04380_ sky130_fd_sc_hd__and2b_1
XANTENNA__11851__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07534_ team_02_WB.instance_to_wrap.top.a1.row2\[15\] net940 _03425_ vssd1 vssd1
+ vccd1 vccd1 _02748_ sky130_fd_sc_hd__o21a_1
XANTENNA__09664__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1 _03405_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout332_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\] net734 net707 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09416__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16810__1364 vssd1 vssd1 vccd1 vccd1 _16810__1364/HI net1364 sky130_fd_sc_hd__conb_1
X_09135_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] net863 _04807_ _04816_
+ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] net697 net677 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08461__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ _03904_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__and2_1
XANTENNA__13079__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold640 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11526__A1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold651 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold662 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold673 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold684 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09968_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\] net661 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a22o_1
X_08919_ _04598_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09899_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] net799 net851 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\]
+ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1340 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 team_02_WB.instance_to_wrap.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2749
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net354 net1727 net543 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07524__B team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11861_ net337 net2357 net549 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16015__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ net1071 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
X_10812_ net378 _06459_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14580_ net1038 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11792_ net332 net2664 net557 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13531_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ _03371_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and3_1
XANTENNA__07540__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _06392_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16250_ clknet_leaf_92_wb_clk_i _02688_ _01207_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_13462_ _03331_ _03332_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__nor2_1
X_10674_ _06325_ _04388_ _04434_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__and3b_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09407__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input95_A wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ clknet_leaf_2_wb_clk_i _01652_ _00159_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12413_ net303 net2173 net490 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__mux2_1
X_16181_ clknet_leaf_72_wb_clk_i _02627_ _01139_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13393_ team_02_WB.instance_to_wrap.top.a1.row1\[15\] _03217_ _03221_ _03226_ team_02_WB.instance_to_wrap.top.a1.row1\[63\]
+ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a32o_1
XANTENNA__12592__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15132_ clknet_leaf_48_wb_clk_i _01583_ _00090_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12962__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ net281 net2180 net498 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ clknet_leaf_84_wb_clk_i _01514_ _00026_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12275_ net266 net2182 net506 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10406__A _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11517__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12714__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ net1022 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
X_11226_ _06736_ _06848_ net383 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XANTENNA__09186__A2 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11936__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _06261_ _06290_ _06292_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ _05760_ _05762_ _05764_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__or4_1
X_15965_ clknet_leaf_117_wb_clk_i _02416_ _00923_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11088_ net428 _06703_ _06720_ _06702_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[21\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14916_ net1162 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
X_10039_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[7\] vssd1 vssd1 vccd1
+ vccd1 _05699_ sky130_fd_sc_hd__or2_1
XANTENNA__11150__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ clknet_leaf_122_wb_clk_i _02347_ _00854_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09894__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ net1155 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11671__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16508__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778_ net1177 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09110__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16517_ clknet_leaf_129_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[20\]
+ _01391_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ net1103 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16448_ clknet_leaf_82_wb_clk_i net2235 _01322_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15532__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16379_ clknet_leaf_73_wb_clk_i _02810_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09377__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12007__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__C_N team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09177__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_61_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout416 net419 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_2
X_09822_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] net675 net635 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a22o_1
XANTENNA__11846__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout427 _06140_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_2
XANTENNA__08924__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ _05413_ _05415_ _05417_ _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__or4_4
XANTENNA__16038__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net747 _04454_ _04466_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09684_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\] net853 net809 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\]
+ _05338_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09885__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08635_ _04402_ _04430_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nor2_1
XANTENNA__10986__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1191_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net914 vssd1 vssd1 vccd1
+ vccd1 _04363_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07517_ net2094 net991 net3 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08497_ _02863_ _04326_ _04279_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout714_A _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08860__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09118_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\] net710 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[28\]
+ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ _04932_ _04951_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09049_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[30\] net823 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09168__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net330 net1919 net530 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
Xhold470 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11756__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _06065_ _06082_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__nand2_1
Xhold492 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__B _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout950 _04553_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout961 _04272_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
Xfanout972 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1 vccd1
+ vccd1 net972 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13121__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _06516_ net226 net942 _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__o211a_1
X_15750_ clknet_leaf_13_wb_clk_i _02201_ _00708_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15405__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A wbm_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ net1167 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
Xhold1181 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ net297 net2570 net540 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XANTENNA__09340__A2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1192 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12587__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ clknet_leaf_0_wb_clk_i _02132_ _00639_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12893_ team_02_WB.instance_to_wrap.top.pc\[4\] _05843_ vssd1 vssd1 vccd1 vccd1 _02927_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ net1158 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11844_ net271 net2506 net551 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
XANTENNA__09628__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14563_ net1068 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15555__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ net263 net1728 net559 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16302_ clknet_leaf_92_wb_clk_i _02735_ _01245_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13514_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] net1690
+ net884 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__o21ai_1
X_10726_ _04972_ net367 vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ net1019 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16233_ clknet_leaf_78_wb_clk_i _00005_ _01190_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13445_ net1650 _03320_ net994 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__o21ai_1
X_10657_ _06232_ _06308_ _06233_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16164_ clknet_leaf_38_wb_clk_i net1621 _01122_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dfrtp_1
X_13376_ net2478 net895 _03278_ net992 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__o211a_1
X_10588_ team_02_WB.instance_to_wrap.top.pc\[25\] _06238_ vssd1 vssd1 vccd1 vccd1
+ _06240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09800__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12327_ net338 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\] net502 vssd1
+ vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__mux2_1
X_15115_ clknet_leaf_20_wb_clk_i _01566_ _00073_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16095_ clknet_leaf_92_wb_clk_i _02541_ _01053_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14831__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ net1161 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09159__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ net326 net2014 net510 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XANTENNA__11666__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11209_ net444 _06830_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12189_ net307 net1788 net519 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
XANTENNA__10174__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ clknet_leaf_22_wb_clk_i _02399_ _00906_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09331__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14278__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15879_ clknet_leaf_16_wb_clk_i _02330_ _00837_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_08420_ team_02_WB.instance_to_wrap.top.a1.row1\[13\] _04285_ vssd1 vssd1 vccd1 vccd1
+ _02714_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10229__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ _04216_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ _04158_ _04160_ _04145_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11441__A3 _06658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_93_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14741__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout497_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout224 _04060_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1204_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
Xfanout246 _06479_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15428__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09570__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _06553_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] net795 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\]
+ _05466_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__a221o_1
Xfanout268 _06891_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
X_07997_ _03845_ _03883_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__xnor2_1
Xfanout279 _06699_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout664_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\] net724 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09322__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _05329_ _05331_ _05333_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15578__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08618_ net977 net931 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__and2b_1
XANTENNA__12200__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _05264_ _05266_ _05267_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08549_ net74 net1612 net892 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11968__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11560_ net351 net2593 net582 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ _05768_ _05791_ _06163_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ _06329_ _07090_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__or2_1
XANTENNA__08633__B _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13230_ net2650 net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[3\]
+ sky130_fd_sc_hd__and2_1
X_10442_ _05543_ net372 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__nand2_1
XANTENNA__09389__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ team_02_WB.instance_to_wrap.top.lcd.currentState\[2\] net985 net896 vssd1
+ vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
X_10373_ _05400_ _06025_ _05357_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12112_ net282 net2089 net588 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input58_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ net230 _03100_ net227 _07052_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__o2bb2a_1
X_12043_ net263 net1716 net531 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10156__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16353__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 _04670_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout791 net792 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15802_ clknet_leaf_121_wb_clk_i _02253_ _00760_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16782_ net1336 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
XANTENNA__09849__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ net1050 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09313__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ clknet_leaf_116_wb_clk_i _02184_ _00691_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ team_02_WB.instance_to_wrap.top.pc\[31\] net946 _07365_ _02978_ vssd1 vssd1
+ vccd1 vccd1 _01529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11120__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12110__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15664_ clknet_leaf_38_wb_clk_i _02115_ _00622_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12876_ team_02_WB.instance_to_wrap.top.pc\[12\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _02910_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14615_ net1156 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11827_ net338 net2571 net554 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15595_ clknet_leaf_21_wb_clk_i _02046_ _00553_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14826__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11758_ net328 net2249 net561 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14546_ net1081 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16689__1243 vssd1 vssd1 vccd1 vccd1 _16689__1243/HI net1243 sky130_fd_sc_hd__conb_1
XFILLER_0_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10709_ _05337_ net374 vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11689_ net310 net2729 net571 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14477_ net1134 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ clknet_leaf_7_wb_clk_i _02661_ _01173_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13428_ net992 _03299_ _03311_ _03309_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13359_ net2624 net895 _03262_ net992 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__o211a_1
X_16147_ clknet_leaf_28_wb_clk_i net1537 _01105_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16078_ clknet_leaf_40_wb_clk_i _02529_ _01036_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07920_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] _03726_ _03764_ vssd1 vssd1
+ vccd1 vccd1 _03811_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ net1189 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__inv_2
XANTENNA__10147__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07851_ _03701_ _03733_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09552__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07563__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07782_ _03637_ _03645_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__and2_1
Xinput2 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_1
X_09521_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[19\] net593 vssd1
+ vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09304__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11111__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09452_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\] net732 net680 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a221o_1
XANTENNA__12020__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08403_ net990 _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09383_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] net801 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout245_A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08334_ _04193_ _04197_ _04210_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16226__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] _04091_ vssd1 vssd1 vccd1
+ vccd1 _04146_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1154_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14471__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09791__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout781_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12703__B _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1010 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_4
Xfanout1019 net1032 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\] net866 net778 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a221o_1
X_10991_ net434 net448 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__nand2_2
XFILLER_0_74_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ _07354_ _07356_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10310__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12661_ _06000_ _06017_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11612_ net296 net2343 net576 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
X_14400_ net1072 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15380_ clknet_leaf_51_wb_clk_i _01831_ _00338_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12592_ net346 net1827 net473 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11810__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ net1048 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ net380 _07095_ _07137_ net386 vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07490__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ net1081 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
X_11474_ net339 net2054 net584 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ team_02_WB.START_ADDR_VAL_REG\[21\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net205 sky130_fd_sc_hd__a21o_1
X_16001_ clknet_leaf_1_wb_clk_i _02452_ _00959_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _04845_ net368 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14193_ net1029 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ _03133_ _03134_ _03135_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__or4_4
XFILLER_0_46_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _05768_ _05792_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__and2_1
XANTENNA__09782__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13075_ net889 _07433_ _03087_ _06993_ net227 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__o32a_1
XANTENNA__12105__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10129__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\] net849 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a22o_1
X_12026_ net326 net1777 net469 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
XANTENNA__09534__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07545__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11944__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15893__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16765_ net1319 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
XFILLER_0_73_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13977_ net1061 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
XANTENNA__13094__A2 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15716_ clknet_leaf_53_wb_clk_i _02167_ _00674_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12928_ _02961_ _02893_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2b_1
X_16696_ net1250 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15647_ clknet_leaf_27_wb_clk_i _02098_ _00605_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12859_ team_02_WB.instance_to_wrap.top.pc\[22\] _06248_ vssd1 vssd1 vccd1 vccd1
+ _02893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15578_ clknet_leaf_116_wb_clk_i _02029_ _00536_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14529_ net1101 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__A0 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _03932_ _03933_ _03907_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a21boi_1
XANTENNA__15273__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10080__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__and2_2
XANTENNA__10324__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ _03787_ _03793_ _03786_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__o21a_1
XANTENNA__09525__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] net915 vssd1 vssd1 vccd1
+ vccd1 _04571_ sky130_fd_sc_hd__or2_1
XANTENNA__08733__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] _03717_ _03718_ vssd1 vssd1
+ vccd1 vccd1 _03725_ sky130_fd_sc_hd__and3_1
XANTENNA__13635__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07765_ _03614_ net350 _03619_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11155__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09504_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\] net868 net799 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
X_07696_ _03542_ _03543_ net362 vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\] net753 _05095_ _05109_
+ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14466__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12045__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _05035_ _05037_ _05039_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or4_2
XFILLER_0_35_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08317_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] net810 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09994__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _04114_ _04116_ _04128_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__or3_2
XANTENNA__10071__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08179_ _04041_ _04062_ _04042_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12899__A2 _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] net686 net639 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11190_ _06059_ _06061_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__nand2_1
XANTENNA__09764__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10141_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[4\] net865 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__09516__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11859__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] net859 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a22o_1
X_16688__1242 vssd1 vssd1 vccd1 vccd1 _16688__1242/HI net1242 sky130_fd_sc_hd__conb_1
XANTENNA__11764__S net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ net1018 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
X_14880_ net1163 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13831_ net1152 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XANTENNA__15146__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12284__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ clknet_leaf_28_wb_clk_i net1415 _01423_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ _06342_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__or2_1
X_13762_ net1093 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ clknet_leaf_23_wb_clk_i _01952_ _00459_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12713_ _04512_ _07339_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__and2_1
X_16481_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[16\] _01355_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12595__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ net1080 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15296__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15432_ clknet_leaf_56_wb_clk_i _01883_ _00390_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12644_ _05977_ _06003_ _06010_ _07172_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15363_ clknet_leaf_40_wb_clk_i _01814_ _00321_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ net279 net1945 net472 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10409__A _05296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08255__A2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14314_ net1027 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ net389 _07038_ net399 vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15294_ clknet_leaf_6_wb_clk_i _01745_ _00252_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11939__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11457_ _06393_ _06398_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__nand2_1
X_14245_ net1087 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15000__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ _05257_ net367 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14176_ net1079 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XANTENNA__09755__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _06146_ _06857_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13127_ _04275_ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] _03126_ vssd1 vssd1
+ vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[7\] sky130_fd_sc_hd__mux2_1
X_10339_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\] net815 _05990_ _05992_
+ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09507__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ _07366_ _03073_ team_02_WB.instance_to_wrap.top.pc\[13\] net945 vssd1 vssd1
+ vccd1 vccd1 _01511_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11674__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ net259 net2369 net470 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
X_16817_ net1371 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
XFILLER_0_75_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16071__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] _03440_ vssd1 vssd1 vccd1
+ vccd1 _03441_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16748_ net1302 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15639__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07481_ net972 net1692 net966 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__10825__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16679_ net1233 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12027__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\] net860 _04899_ vssd1
+ vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09151_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\] net638 _04831_ vssd1
+ vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15789__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ _03951_ net225 _03956_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09082_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[29\] net879 net875 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a22o_1
XANTENNA__10053__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11849__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _03877_ _03911_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput60 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
XFILLER_0_115_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold800 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput71 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_1
XFILLER_0_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold811 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold822 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold833 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold844 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold855 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold866 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold877 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold888 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09984_ _05639_ _05641_ _05643_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__or4_1
Xhold899 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1117_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08935_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\] net710 net680 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\]
+ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07509__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16414__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout577_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ net959 _04296_ _04308_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07817_ _03706_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__or2_1
X_08797_ net168 net952 net903 net1560 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout744_A _06323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ _03577_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09131__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07679_ _03560_ _03562_ _03567_ _03565_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08485__A2 _04315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09418_ _05086_ _05088_ _05090_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__or4_1
X_10690_ team_02_WB.instance_to_wrap.top.pc\[25\] team_02_WB.instance_to_wrap.top.pc\[24\]
+ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09349_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] net871 net799 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ net337 net2685 net498 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__mux2_1
XANTENNA__10044__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11759__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ net435 _06920_ _06927_ net440 _06925_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__o221a_1
X_12291_ net327 net2661 net505 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08641__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14030_ net1063 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07538__A team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11242_ _06178_ _06862_ _06149_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09737__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ net437 _06799_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input40_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\] net807 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a22o_1
X_15981_ clknet_leaf_33_wb_clk_i _02432_ _00939_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13297__A2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10055_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] net693 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__a22o_1
X_14932_ net1001 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__09370__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ net1172 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ clknet_leaf_61_wb_clk_i _02836_ _01475_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ net1109 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14794_ net1174 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16533_ clknet_leaf_129_wb_clk_i net1403 _01406_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ net1030 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ _06079_ _06081_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__nand2_1
XANTENNA__08476__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16464_ clknet_leaf_67_wb_clk_i net1487 _01338_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10283__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13676_ net1005 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10888_ _04804_ net373 _06078_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__a21bo_1
X_15415_ clknet_leaf_116_wb_clk_i _01866_ _00373_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12627_ net410 _06811_ _06813_ _06799_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__o211a_1
X_16395_ clknet_leaf_74_wb_clk_i _02826_ _01269_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10035__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ clknet_leaf_25_wb_clk_i _01797_ _00304_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09976__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12558_ net339 net2416 net464 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11669__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ _06161_ _07107_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ clknet_leaf_23_wb_clk_i _01728_ _00235_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__B _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12489_ net328 net2112 net481 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__mux2_1
Xhold107 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\] vssd1 vssd1 vccd1 vccd1
+ net1505 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[3\] vssd1 vssd1 vccd1
+ vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold129 _02607_ vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14228_ net1052 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XANTENNA__09728__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08936__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15311__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14159_ net1126 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08400__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13288__A2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ net1465 net988 _04438_ _04516_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12496__A0 _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09361__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1184 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_2
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_4
X_08651_ net746 _04445_ _04446_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09900__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _03461_ _03490_ _03463_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net973 net975 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07533_ net2618 net935 net918 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ net6 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] net738 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout325_A _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1067_A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\] net806 net786 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16687__1241 vssd1 vssd1 vccd1 vccd1 _16687__1241/HI net1241 sky130_fd_sc_hd__conb_1
XANTENNA__10026__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09838__A _05493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09967__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10991__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[29\] net721 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\]
+ _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08016_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _03869_ net241 vssd1 vssd1
+ vccd1 vccd1 _03905_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09719__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold630 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold652 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] vssd1 vssd1 vccd1 vccd1
+ net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold685 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold696 team_02_WB.instance_to_wrap.top.pad.keyCode\[2\] vssd1 vssd1 vccd1 vccd1
+ net2094 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15804__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] net702 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\]
+ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout861_A _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _04601_ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__nand2_2
XANTENNA__12203__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] net871 net807 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a22o_1
Xhold1330 team_02_WB.instance_to_wrap.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net2728
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09352__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1352 team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net2750
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ net38 net947 net921 net2681 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ net335 net2274 net548 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XANTENNA__09104__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11791_ net327 net2565 net557 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13530_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] _03373_
+ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__or2_1
XANTENNA__07540__B team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10265__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10742_ _05677_ net375 vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ net826 net581 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nand2_1
X_13461_ net1684 _03330_ net994 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ clknet_leaf_10_wb_clk_i _01651_ _00158_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12412_ net297 net2387 net488 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__mux2_1
X_16180_ clknet_leaf_71_wb_clk_i _02626_ _01138_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11214__B2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input88_A wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13392_ _03274_ _03289_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15131_ clknet_leaf_119_wb_clk_i _01582_ _00089_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15334__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ net274 net2328 net499 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ net261 net2002 net507 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__mux2_1
X_15062_ clknet_leaf_81_wb_clk_i _01513_ _00025_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12714__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11517__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ _06789_ _06847_ net377 vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__mux2_1
X_14013_ net1055 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09591__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11156_ _06257_ net744 net458 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _06782_
+ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\] net686 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\]
+ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a221o_1
X_15964_ clknet_leaf_63_wb_clk_i _02415_ _00922_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11087_ net409 net450 _06713_ _06719_ _06707_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a311o_1
XANTENNA__10422__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12113__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ net1158 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_10038_ _05690_ _05694_ _05696_ _05698_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[7\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_136_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15895_ clknet_leaf_120_wb_clk_i _02346_ _00853_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08697__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14846_ net1155 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16466__D team_02_WB.instance_to_wrap.top.aluOut\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14777_ net1179 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
X_11989_ net1920 net301 net534 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16516_ clknet_leaf_28_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[19\]
+ _01390_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10256__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13728_ net1070 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16447_ clknet_leaf_81_wb_clk_i net1466 _01321_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13659_ net1047 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14564__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16378_ clknet_leaf_73_wb_clk_i _02809_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15329_ clknet_leaf_1_wb_clk_i _01780_ _00287_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15827__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_2
X_09821_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\] net659 net651 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a221o_1
XANTENNA__09582__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_2
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
Xfanout439 _06056_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15977__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09752_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\] net636 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a221o_1
XANTENNA__12023__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ net747 _04449_ _04466_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09683_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\] net845 _05350_ _05351_
+ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a211o_1
XANTENNA__08688__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08634_ _04394_ _04395_ _04396_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15207__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08565_ team_02_WB.instance_to_wrap.top.a1.instruction\[3\] net914 vssd1 vssd1 vccd1
+ vccd1 _04362_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout442_A _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ net1959 net991 net4 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a21o_1
XANTENNA__10247__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08496_ net2713 _04331_ _04325_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16602__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_A _04461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12944__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09117_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] net721 net694 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[30\] net870 net802 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\]
+ _04724_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold460 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12722__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold482 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _06040_ _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__xnor2_1
Xhold493 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10183__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 _03421_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_2
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout962 net971 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_2
Xfanout984 team_02_WB.instance_to_wrap.top.ru.dmmRen vssd1 vssd1 vccd1 vccd1 net984
+ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 _00012_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09325__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12961_ _07370_ _07371_ _02868_ _02869_ net888 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08679__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net1163 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ net289 net1847 net540 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
X_15680_ clknet_leaf_6_wb_clk_i _02131_ _00638_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1193 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ _02924_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ net1158 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net276 net2541 net550 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14562_ net1090 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11774_ net261 net1979 net558 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16301_ clknet_leaf_90_wb_clk_i _02734_ _01244_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13513_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\] net884
+ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10725_ _05012_ net375 vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14493_ net1055 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
XANTENNA__08851__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16232_ clknet_leaf_28_wb_clk_i _00010_ _01189_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dfrtp_2
X_13444_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\] _03320_ vssd1 vssd1 vccd1
+ vccd1 _03321_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10656_ team_02_WB.instance_to_wrap.top.pc\[26\] _06235_ _06307_ vssd1 vssd1 vccd1
+ vccd1 _06308_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ clknet_leaf_28_wb_clk_i net1657 _01121_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dfrtp_1
X_10587_ team_02_WB.instance_to_wrap.top.pc\[25\] _06238_ vssd1 vssd1 vccd1 vccd1
+ _06239_ sky130_fd_sc_hd__or2_1
XANTENNA__12108__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13375_ _03264_ _03270_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__or3b_1
XFILLER_0_134_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15114_ clknet_leaf_44_wb_clk_i _01565_ _00072_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12326_ _07055_ net1883 net501 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
X_16094_ clknet_leaf_92_wb_clk_i _02540_ _01052_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11947__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ net1162 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__inv_2
X_12257_ net313 net2218 net510 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11208_ _06290_ _06831_ net909 vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3b_1
X_12188_ net299 net1782 net518 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _05196_ net431 _06583_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13112__A1 _07410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15947_ clknet_leaf_20_wb_clk_i _02398_ _00905_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16686__1240 vssd1 vssd1 vccd1 vccd1 _16686__1240/HI net1240 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15878_ clknet_leaf_15_wb_clk_i _02329_ _00836_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14829_ net1190 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16625__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ _04209_ _04215_ _04201_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ _04158_ _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08842__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13402__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11857__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07566__C1 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 _03968_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout392_A _05908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11362__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _07186_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
Xfanout247 _06479_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_1
X_09804_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] net803 net766 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\]
+ _05465_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a221o_1
Xfanout258 net261 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout269 _06891_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ _03884_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nor2_1
XANTENNA__16155__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ _05399_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__and2b_1
XANTENNA__11114__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13373__A _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09666_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\] net712 net680 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\]
+ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08617_ _04389_ _04390_ _04408_ _04375_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09597_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] net803 net844 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ _05258_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout824_A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ net75 net1644 net891 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XANTENNA__09086__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08479_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.row1\[111\]
+ net752 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XANTENNA__08833__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12717__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire604 _05611_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_2
X_10510_ _05768_ _05791_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11490_ team_02_WB.instance_to_wrap.top.pc\[5\] _06328_ vssd1 vssd1 vccd1 vccd1 _07090_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ _05503_ net367 vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__nand2_1
XANTENNA__08046__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13160_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] team_02_WB.instance_to_wrap.top.lcd.currentState\[0\]
+ _03137_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
X_10372_ _05402_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net273 net1735 net588 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XANTENNA__11767__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13091_ _07406_ _07425_ _07427_ net890 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__o31ai_1
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09546__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net259 net1957 net529 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
Xhold290 net141 vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09010__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 _04673_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
X_15801_ clknet_leaf_112_wb_clk_i _02252_ _00759_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout781 _04669_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_8
Xfanout792 _04663_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16781_ net1335 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13993_ net1024 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XANTENNA__15522__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ clknet_leaf_54_wb_clk_i _02183_ _00690_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ net231 _02976_ _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10700__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15663_ clknet_leaf_31_wb_clk_i _02114_ _00621_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12875_ _02907_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nand2_1
X_14614_ net1158 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11826_ net334 net2532 net552 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15594_ clknet_leaf_51_wb_clk_i _02045_ _00552_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09077__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14545_ net1078 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11757_ net312 net2457 net561 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08824__B net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10092__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ _06357_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14476_ net1019 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
X_11688_ net301 net2113 net569 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16215_ clknet_leaf_36_wb_clk_i _02660_ _01172_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13427_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__or2_1
X_10639_ team_02_WB.instance_to_wrap.top.pc\[18\] _06257_ vssd1 vssd1 vccd1 vccd1
+ _06291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16146_ clknet_leaf_6_wb_clk_i net1534 _01104_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13358_ _03254_ _03257_ _03261_ _03210_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__or4b_2
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11677__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ net275 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\] net500 vssd1
+ vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__mux2_1
X_16077_ clknet_leaf_33_wb_clk_i _02528_ _01035_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13289_ _03181_ _03185_ _03179_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15052__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09537__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15028_ net1164 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09001__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07850_ _03709_ _03736_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_120_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ _03660_ _03667_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__nand2_1
Xinput3 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
X_09520_ _05186_ _05190_ _05191_ _05192_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[19\]
+ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\] net708 net692 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08402_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03417_ vssd1 vssd1 vccd1
+ vccd1 _04269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09382_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] net869 net841 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a22o_1
XANTENNA__09068__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08333_ _04189_ _04196_ _04191_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__o21a_1
XANTENNA__08815__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ _04134_ _04137_ _04143_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ _04077_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1147_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09528__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08751__B2 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _03867_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09718_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\] net846 net875 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a22o_1
XANTENNA__12211__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ net408 _06626_ _06628_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_39_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _05316_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__and2b_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12660_ _05570_ _06127_ _07285_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__or4_1
XANTENNA_input105_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ net289 net2361 net576 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12591_ net337 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\] net473 vssd1
+ vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08806__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ net1046 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
XANTENNA__10074__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11542_ net380 _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ net1117 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11473_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[6\] _07074_ vssd1 vssd1 vccd1
+ vccd1 _07075_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15075__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16000_ clknet_leaf_8_wb_clk_i _02451_ _00958_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13212_ team_02_WB.START_ADDR_VAL_REG\[20\] _04356_ vssd1 vssd1 vccd1 vccd1 net204
+ sky130_fd_sc_hd__and2_1
XANTENNA_input70_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09767__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ net378 _06074_ _06075_ _06076_ net384 vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ net1016 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or4b_1
X_10355_ _05884_ _06007_ _05839_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13074_ _07402_ _07432_ _07401_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__a21oi_1
X_10286_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\] net865 net797 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\]
+ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12025_ net312 net2166 net469 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
XANTENNA__16470__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A2 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16764_ net1318 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
XANTENNA__12121__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ net1107 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
XANTENNA__09298__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ clknet_leaf_45_wb_clk_i _02166_ _00673_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12927_ _02896_ _02897_ _02959_ _02894_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a31o_1
X_16695_ net1249 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__10301__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11960__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13741__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15646_ clknet_leaf_6_wb_clk_i _02097_ _00604_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12858_ team_02_WB.instance_to_wrap.top.pc\[22\] _06248_ vssd1 vssd1 vccd1 vccd1
+ _02892_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ net275 net2537 net553 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15577_ clknet_leaf_107_wb_clk_i _02028_ _00535_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12789_ _07337_ _07341_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15418__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528_ net1075 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09470__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14459_ net1060 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09758__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15568__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ clknet_leaf_66_wb_clk_i _02575_ _01087_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] _04635_ vssd1 vssd1
+ vccd1 vccd1 _04636_ sky130_fd_sc_hd__and2b_2
XANTENNA__10324__B _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07902_ _03790_ _03791_ _03783_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21o_1
X_08882_ net1562 _04570_ net825 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08733__B2 _04523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _03717_ _03718_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1
+ vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12031__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _03614_ _03619_ net350 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09289__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\] net881 net877 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07695_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _03582_ _03583_ _03584_ vssd1
+ vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout355_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14747__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] net805 net793 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\]
+ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] net722 net670 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\]
+ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_A _07212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15098__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08316_ _04178_ _04184_ _04187_ _04192_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\] net813 net786 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08247_ _04116_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09749__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _04058_ net224 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09213__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12206__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\] net880 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[25] sky130_fd_sc_hd__clkbuf_4
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
X_10071_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] net811 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09921__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ net1092 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
XANTENNA__07543__B team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11087__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ net1146 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
X_10973_ team_02_WB.instance_to_wrap.top.pc\[24\] _06341_ team_02_WB.instance_to_wrap.top.pc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11780__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15500_ clknet_leaf_52_wb_clk_i _01951_ _00458_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10295__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _04512_ _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16480_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[15\] _01354_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13692_ net1097 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ clknet_leaf_114_wb_clk_i _01882_ _00389_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _06154_ _07239_ _07265_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10047__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ clknet_leaf_47_wb_clk_i _01813_ _00320_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12574_ net272 net2245 net474 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09452__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ net1012 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ net376 _07080_ _07121_ net383 vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__o211a_1
XANTENNA__15710__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15293_ clknet_leaf_111_wb_clk_i _01744_ _00251_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ net1143 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11456_ _06013_ _07058_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__nor2_1
XANTENNA__09204__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _06058_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12116__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14175_ net1130 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
X_11387_ net313 net2325 net584 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XANTENNA__10425__A _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ net1667 _03126_ _03128_ net990 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15860__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10338_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\] net779 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__S net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13057_ _06931_ net227 _03072_ net889 _03070_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o221a_1
X_10269_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[2\] net680 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07518__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ net254 net2435 net470 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XANTENNA__09912__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16216__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16816_ net1370 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
X_13959_ net1153 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
X_16747_ net1301 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14567__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11690__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07480_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] team_02_WB.instance_to_wrap.ramload\[25\]
+ net964 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
X_16678_ net1232 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__15240__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__A team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16366__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15629_ clknet_leaf_23_wb_clk_i _02080_ _00587_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09150_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\] net634 net619 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a22o_1
XANTENNA__09979__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09443__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__inv_2
XANTENNA__15390__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13410__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08032_ _03876_ _03911_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput61 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
Xhold801 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput72 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
Xhold812 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput83 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold823 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput94 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12026__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold867 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold878 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold889 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\] net799 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a221o_1
XANTENNA__11865__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] net724 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1012_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08865_ net1578 _04560_ net825 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__mux2_1
XANTENNA__10513__A1 _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ _03667_ _03694_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08796_ net169 net952 net903 net1553 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
X_07747_ _03580_ _03601_ _03604_ _03581_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a22o_1
XANTENNA__14477__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07678_ _03560_ net362 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09682__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12709__B _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] net696 net692 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\]
+ _05091_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a221o_1
XANTENNA__13215__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15733__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\] net775 net760 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09434__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09279_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\] net645 net617 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a221o_1
X_11310_ _06149_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12290_ net313 net2450 net505 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11241_ _05484_ _06861_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__or2_1
XANTENNA__07538__B team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10201__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11172_ _06797_ _06798_ net410 vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _05776_ _05778_ _05780_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or4_1
X_15980_ clknet_leaf_53_wb_clk_i _02431_ _00938_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13151__C1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A wbm_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ net1042 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XANTENNA__07554__A team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10054_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] net714 net661 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\]
+ _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a221o_1
X_14862_ net1173 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13813_ net1120 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_16601_ clknet_leaf_75_wb_clk_i _02835_ _01474_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_14793_ net1174 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10268__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16532_ clknet_leaf_7_wb_clk_i net1457 _01405_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13744_ net1017 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
X_10956_ net408 _06596_ _06593_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08385__A team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16463_ clknet_leaf_65_wb_clk_i net1701 _01337_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13675_ net1014 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
X_10887_ net408 _06530_ _06527_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15414_ clknet_leaf_110_wb_clk_i _01865_ _00372_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12626_ _06661_ _06688_ _06734_ _06706_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__or4b_1
X_16394_ clknet_leaf_74_wb_clk_i _02825_ _01268_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09425__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15345_ clknet_leaf_17_wb_clk_i _01796_ _00303_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12557_ net335 net2607 net465 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _05839_ _06160_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__nand2_1
X_15276_ clknet_leaf_52_wb_clk_i _01727_ _00234_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ net311 net2530 net482 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold108 team_02_WB.instance_to_wrap.top.pc\[13\] vssd1 vssd1 vccd1 vccd1 net1506
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 _02582_ vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ net1148 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11439_ net417 _06652_ _07042_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13390__C1 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14158_ net1065 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11685__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ team_02_WB.instance_to_wrap.top.pc\[4\] net945 net941 _03115_ vssd1 vssd1
+ vccd1 vccd1 _01502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14089_ net1012 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07464__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1170 net1205 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ net747 _04445_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__and3_4
XFILLER_0_59_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1181 net1183 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_4
Xfanout1192 net1204 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__buf_2
X_07601_ _03441_ _03484_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08581_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_87_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15756__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10259__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13405__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07532_ _03419_ net940 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09664__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ net1175 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09202_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] net730 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11759__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09416__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09133_ _04810_ _04811_ _04813_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09838__B _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09064_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] net662 net645 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15136__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08461__C _04315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08015_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] net241 _03869_ vssd1 vssd1
+ vccd1 vccd1 _03904_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold620 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold642 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold653 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\] vssd1
+ vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold686 team_02_WB.instance_to_wrap.top.pad.keyCode\[6\] vssd1 vssd1 vccd1 vccd1
+ net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold697 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\] net738 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08917_ _04392_ _04594_ _04384_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__o21ai_4
XANTENNA__16531__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\] net822 net855 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\]
+ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a221o_1
Xhold1320 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout854_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1331 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ net8 net949 net923 net2065 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
Xhold1342 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08779_ net1679 net956 net927 _04546_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
X_10810_ _04722_ net368 _06073_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11790_ net313 net2644 net556 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09655__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ _05633_ net370 vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10670__B1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] _03330_ vssd1 vssd1 vccd1
+ vccd1 _03331_ sky130_fd_sc_hd__and2_1
X_10672_ _04388_ net826 _04434_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09407__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ net288 net2072 net488 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13391_ net1566 net895 _03290_ net992 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08652__B team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15130_ clknet_leaf_120_wb_clk_i _01581_ _00088_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12962__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ net277 net2277 net497 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10973__A1 team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16061__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15061_ clknet_leaf_84_wb_clk_i _01512_ _00024_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_12273_ net255 net2040 net506 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15629__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14012_ net1084 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
X_11224_ _06357_ _06361_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09040__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11155_ net911 _06781_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nor2_1
XANTENNA__10703__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[5\] net722 net705 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15963_ clknet_leaf_118_wb_clk_i _02414_ _00921_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11086_ _06034_ net433 _06580_ _06717_ _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10422__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15779__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14914_ net1150 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
X_10037_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] net789 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\]
+ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a221o_1
X_15894_ clknet_leaf_111_wb_clk_i _02345_ _00852_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14845_ net1155 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15006__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14776_ net1181 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
X_11988_ net2306 net291 net532 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09646__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16515_ clknet_leaf_38_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[18\]
+ _01389_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13727_ net1125 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08854__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ net445 _06581_ _04912_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13658_ net1052 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
X_16446_ clknet_leaf_81_wb_clk_i net1506 _01320_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ _06440_ _06523_ _07236_ _06481_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__or4b_1
X_16377_ clknet_leaf_73_wb_clk_i _02808_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16482__D team_02_WB.instance_to_wrap.top.aluOut\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13589_ net1161 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15328_ clknet_leaf_8_wb_clk_i _01779_ _00286_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15259_ clknet_leaf_119_wb_clk_i _01710_ _00217_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16554__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] net711 net639 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a22o_1
Xfanout407 _05862_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12304__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout429 _06139_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10192__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09751_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\] net708 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__a22o_1
X_08702_ net745 _04446_ _04466_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and3_1
X_09682_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\] net874 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[15\]
+ _05340_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__a221o_1
XANTENNA__09885__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _04367_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout268_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ net979 _04359_ net977 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07515_ net2329 net116 _00011_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08845__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04269_ _04274_ _04279_
+ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__o311a_1
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1177_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09116_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] net662 net645 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\]
+ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09270__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\] net878 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\]
+ _04727_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09022__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold483 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12214__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold494 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15921__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779__1333 vssd1 vssd1 vccd1 vccd1 _16779__1333/HI net1333 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
X_09949_ net604 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[9\]
+ sky130_fd_sc_hd__inv_2
Xfanout952 net954 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net971 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_2
Xfanout974 team_02_WB.instance_to_wrap.top.a1.instruction\[14\] vssd1 vssd1 vccd1
+ vccd1 net974 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1
+ net985 sky130_fd_sc_hd__buf_2
XANTENNA__13121__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12960_ net229 _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nand2_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1150 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09876__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1161 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ net280 net1789 net540 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ team_02_WB.instance_to_wrap.top.pc\[5\] _05797_ vssd1 vssd1 vccd1 vccd1 _02925_
+ sky130_fd_sc_hd__or2_1
Xhold1183 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 team_02_WB.instance_to_wrap.top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 net2592
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ net1156 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11842_ net265 net1841 net550 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09089__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14561_ net1102 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08836__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ net254 net1762 net558 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XANTENNA__15301__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16427__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13512_ _03361_ _03362_ _03363_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__and3_1
X_16300_ clknet_leaf_98_wb_clk_i _02733_ _01243_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ _06373_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__nand2_1
X_16735__1289 vssd1 vssd1 vccd1 vccd1 _16735__1289/HI net1289 sky130_fd_sc_hd__conb_1
X_14492_ net1124 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16231_ clknet_leaf_28_wb_clk_i _02676_ _01188_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13443_ net1176 _03319_ _03320_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nor3_1
X_10655_ _06236_ _06239_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16162_ clknet_leaf_38_wb_clk_i net1640 _01120_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ _03206_ _03276_ _03137_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09261__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10586_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net930 net591 vssd1
+ vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09800__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15113_ clknet_leaf_31_wb_clk_i _01564_ _00071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12325_ net332 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\] net502 vssd1
+ vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
X_16093_ clknet_leaf_92_wb_clk_i _02539_ _01051_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15044_ net1162 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__inv_2
X_12256_ net307 net2446 net511 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _06264_ _06287_ _06289_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__or3b_1
XANTENNA__13360__A2 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12124__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ net293 net1774 net516 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XANTENNA__10174__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _05194_ net447 _06184_ net452 vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a22o_1
XANTENNA__11963__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15946_ clknet_leaf_46_wb_clk_i _02397_ _00904_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ net440 _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09867__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16477__D team_02_WB.instance_to_wrap.top.aluOut\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15877_ clknet_leaf_127_wb_clk_i _02328_ _00835_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14828_ net1188 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09619__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08827__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14759_ net1178 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ _04149_ _04152_ _04150_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16429_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[28\]
+ _01303_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15944__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12034__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _07336_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10165__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
X_09803_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\] net787 net775 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a221o_1
XANTENNA__11362__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _06479_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ _03845_ _03883_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout385_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _05378_ _05397_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09665_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] net696 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a22o_1
XANTENNA__15324__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08616_ net977 net910 _04411_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__and4_1
X_09596_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] net852 net760 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\]
+ _05262_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08547_ net76 team_02_WB.START_ADDR_VAL_REG\[13\] net894 vssd1 vssd1 vccd1 vccd1
+ _02658_ sky130_fd_sc_hd__mux2_1
XANTENNA__08818__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout817_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08478_ net1615 net751 net742 _04297_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
XANTENNA__09491__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12209__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08046__A1 team_02_WB.instance_to_wrap.top.a1.row2\[41\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _06089_ _06092_ net363 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _06021_ _06023_ _05441_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ net276 net2150 net587 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13090_ _02920_ _02937_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12041_ net256 net2373 net531 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
Xhold280 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_02_WB.instance_to_wrap.ramload\[21\] vssd1 vssd1 vccd1 vccd1 net1689
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10156__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11783__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _04679_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15800_ clknet_leaf_121_wb_clk_i _02251_ _00758_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13564__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 _04673_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_6
Xfanout782 _04669_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16780_ net1334 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
X_13992_ net1099 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
Xfanout793 _04661_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_6
XFILLER_0_137_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09849__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12943_ _06346_ net226 _02875_ _04363_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o22a_1
X_15731_ clknet_leaf_125_wb_clk_i _02182_ _00689_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10700__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11084__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15662_ clknet_leaf_40_wb_clk_i _02113_ _00620_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12874_ team_02_WB.instance_to_wrap.top.pc\[13\] _06276_ vssd1 vssd1 vccd1 vccd1
+ _02908_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15817__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613_ net1156 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11825_ net332 net2498 net554 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
XANTENNA__08809__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15593_ clknet_leaf_24_wb_clk_i _02044_ _00551_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ net1018 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
X_11756_ net309 net2517 net562 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07501__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _05215_ net368 vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__nand2_1
X_14475_ net1027 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XANTENNA__10428__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ net293 net2104 net568 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__mux2_1
XANTENNA__12119__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16214_ clknet_leaf_36_wb_clk_i _02659_ _01171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13426_ net1597 _03310_ net1176 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a21oi_1
X_10638_ _06264_ _06287_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ clknet_leaf_0_wb_clk_i net1520 _01103_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11958__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ team_02_WB.instance_to_wrap.top.a1.row1\[106\] _03216_ _03258_ _03260_ vssd1
+ vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ net928 _04629_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and2b_1
XANTENNA__11592__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ net265 net2004 net503 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16076_ clknet_leaf_52_wb_clk_i _02527_ _01034_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13288_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\] _03174_ _03187_ _03198_
+ net995 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15027_ net1154 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ net251 net1936 net509 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10147__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09952__A _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15347__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07780_ _03631_ _03666_ _03667_ _03669_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_21_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15929_ clknet_leaf_117_wb_clk_i _02380_ _00887_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ _05117_ _05119_ _05121_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__or4_2
XFILLER_0_137_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08401_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09381_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] net862 net807 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09399__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _04185_ _04202_ _04203_ _04207_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16778__1332 vssd1 vssd1 vccd1 vccd1 _16778__1332/HI net1332 sky130_fd_sc_hd__conb_1
XFILLER_0_34_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08263_ _04137_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12029__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ _04057_ net224 _04045_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09225__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13021__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16122__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16734__1288 vssd1 vssd1 vccd1 vccd1 _16734__1288/HI net1288 sky130_fd_sc_hd__conb_1
XFILLER_0_96_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout767_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13088__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03858_ _03859_ vssd1 vssd1
+ vccd1 vccd1 _03868_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\] net818 net834 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout934_A _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _05296_ _05315_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10310__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] net718 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11610_ net280 net1758 net576 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12590_ net335 net2441 net472 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09464__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09102__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__B1 team_02_WB.instance_to_wrap.top.aluOut\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _05883_ _05929_ net369 vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14260_ net1053 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] net887 net907 team_02_WB.instance_to_wrap.top.pc\[6\]
+ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09216__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ team_02_WB.START_ADDR_VAL_REG\[19\] net998 _04355_ vssd1 vssd1 vccd1 vccd1
+ net202 sky130_fd_sc_hd__a21o_1
XFILLER_0_122_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11778__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _04722_ net368 net378 vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14191_ net1110 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07557__A team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13142_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input63_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10354_ _06002_ _06006_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and2_1
X_13073_ _02942_ _03085_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__xnor2_1
X_10285_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\] net857 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a22o_1
XANTENNA__10129__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ net307 net2735 net471 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12402__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout590 _06221_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ net1317 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
X_13975_ net1108 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
X_15714_ clknet_leaf_49_wb_clk_i _02165_ _00672_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ _02897_ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__nand2_1
X_16694_ net1248 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_38_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10301__A2 _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ clknet_leaf_111_wb_clk_i _02096_ _00603_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ _02889_ _02890_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ net263 net1895 net553 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15576_ clknet_leaf_123_wb_clk_i _02027_ _00534_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09455__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12788_ _07410_ _07411_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14527_ net1132 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11739_ net250 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net562 vssd1
+ vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14458_ net1052 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13003__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11688__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16490__D team_02_WB.instance_to_wrap.top.aluOut\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13409_ net1475 _04228_ net828 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
X_14389_ net1119 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07467__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ clknet_leaf_65_wb_clk_i _02574_ _01086_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08950_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] net886 vssd1 vssd1 vccd1
+ vccd1 _04635_ sky130_fd_sc_hd__and2_1
X_16059_ clknet_leaf_104_wb_clk_i _02510_ _01017_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11317__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08881_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] net939 _04568_ _04569_ vssd1
+ vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13408__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09930__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07763_ _03650_ _03653_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ _05168_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07694_ _03583_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and2_1
XANTENNA__09694__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] net797 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout250_A _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09364_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[22\] net664 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a22o_1
XANTENNA__09446__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08315_ _04189_ _04191_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09295_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] net823 net778 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A _07215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _04107_ _04118_ _04096_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15512__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _04058_ net224 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12753__B1 _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15662__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
X_10070_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] net847 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12222__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ net1071 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
X_10972_ _06239_ _06240_ _06305_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__a21o_1
XANTENNA__09685__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _07337_ _07338_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__nor2_1
X_13691_ net1048 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12642_ _05703_ _05749_ _05839_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__or4_1
X_15430_ clknet_leaf_12_wb_clk_i _01881_ _00388_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ clknet_leaf_130_wb_clk_i _01812_ _00319_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12573_ net275 net2302 net474 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12992__B1 team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11524_ net380 _07120_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__nand2_1
X_14312_ net1089 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
X_15292_ clknet_leaf_63_wb_clk_i _01743_ _00250_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14243_ net1073 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ _05749_ _05793_ _06012_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__nor3_1
XFILLER_0_81_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10706__A _05257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10406_ _05215_ net372 vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14174_ net1020 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ net459 team_02_WB.instance_to_wrap.top.aluOut\[10\] _06995_ _06887_ vssd1
+ vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__o22a_4
XANTENNA__10425__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13125_ _04269_ _03126_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10337_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\] net796 net787 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13056_ _07437_ _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10268_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\] net692 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a22o_1
XANTENNA__08176__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ net250 net2575 net470 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
X_16777__1331 vssd1 vssd1 vccd1 vccd1 _16777__1331/HI net1331 sky130_fd_sc_hd__conb_1
XANTENNA__10441__A _05503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\] net820 _05853_ _05855_
+ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a211o_1
XANTENNA__07923__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16815_ net1369 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
XFILLER_0_89_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11971__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16746_ net1300 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
X_13958_ net1139 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XANTENNA__09676__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12909_ team_02_WB.instance_to_wrap.top.pc\[10\] _05593_ _02942_ vssd1 vssd1 vccd1
+ vccd1 _02943_ sky130_fd_sc_hd__o21a_1
X_16677_ net1231 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_124_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13889_ net1143 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XANTENNA__08565__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15628_ clknet_leaf_52_wb_clk_i _02079_ _00586_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09428__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15559_ clknet_leaf_16_wb_clk_i _02010_ _00517_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16733__1287 vssd1 vssd1 vccd1 vccd1 _16733__1287/HI net1287 sky130_fd_sc_hd__conb_1
X_08100_ _03984_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _04753_ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__nor2_8
XFILLER_0_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08031_ _03880_ _03912_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12307__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput62 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11211__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
XANTENNA__15685__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold824 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09600__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold835 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11214__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13927__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold868 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] net807 net766 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a22o_1
Xhold879 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\] net694 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12042__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net959 _04293_ _04305_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a32o_1
XANTENNA__10351__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1005_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07815_ _03657_ _03705_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__xnor2_2
X_08795_ net170 net953 net904 net1510 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11881__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1113_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07746_ _03614_ _03620_ _03628_ _03633_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09131__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07677_ _03560_ _03566_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout632_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] net724 net716 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] net864 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09278_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] net665 net633 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12725__B _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08229_ _04086_ _04111_ _04090_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12217__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12726__B1 _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _06148_ _06860_ _06171_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11171_ _06570_ _06574_ net404 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__mux2_1
XANTENNA__12741__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10122_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\] net862 net779 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\]
+ _05773_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10053_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\] net734 net722 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a22o_1
X_14930_ net1003 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XANTENNA__15408__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__A2 _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A wbm_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1173 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11791__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ clknet_leaf_82_wb_clk_i _02834_ _01473_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13812_ net1038 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
X_14792_ net1173 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XANTENNA__11465__B1 _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16531_ clknet_leaf_6_wb_clk_i net1435 _01404_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13743_ net1123 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
X_10955_ _06594_ _06595_ net403 vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16462_ clknet_leaf_65_wb_clk_i net1607 _01336_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13674_ net1036 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XANTENNA__08881__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15413_ clknet_leaf_115_wb_clk_i _01864_ _00371_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12625_ _06500_ _06410_ _06118_ _06457_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__or4bb_1
X_16393_ clknet_leaf_77_wb_clk_i _02824_ _01267_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15344_ clknet_leaf_34_wb_clk_i _01795_ _00302_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ net330 net2025 net464 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ net437 _07105_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__nor2_1
X_12487_ net307 net1907 net482 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__mux2_1
X_15275_ clknet_leaf_21_wb_clk_i _01726_ _00233_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12127__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[5\] vssd1 vssd1 vccd1 vccd1
+ net1507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11438_ net417 _06654_ _07042_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a21oi_1
X_14226_ net1084 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11966__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ net1132 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XANTENNA__08936__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11369_ _06940_ _06979_ net380 vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13108_ _07113_ net228 _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__o21ai_1
X_14088_ net1100 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
X_13039_ net888 _07442_ _03056_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09897__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1205 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09361__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1182 net1183 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
Xfanout1193 net1195 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_4
X_07600_ _03461_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13482__A _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08580_ net973 net975 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09113__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07531_ _03418_ net936 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16729_ net1283 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16483__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ team_02_WB.instance_to_wrap.top.edg2.flip2 vssd1 vssd1 vccd1 vccd1 _03403_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_9_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08872__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09201_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\] net670 net643 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09132_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\] net830 net758 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ _04808_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a221o_1
XANTENNA__09821__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09063_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[29\] net737 net653 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\]
+ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a221o_1
XANTENNA__12037__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__A _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] net241 vssd1 vssd1 vccd1 vccd1
+ _03903_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold610 team_02_WB.instance_to_wrap.top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1 net2008
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11876__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold654 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold665 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09965_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\] net650 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\]
+ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout582_A _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net910 _04599_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nand2_1
X_09896_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net791 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a22o_1
XANTENNA__09888__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1310 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 team_02_WB.instance_to_wrap.top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1 net2719
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1332 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09352__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net9 net948 net922 net1713 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__o22a_1
Xhold1343 team_02_WB.instance_to_wrap.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net2741
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout847_A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15700__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13436__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08778_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[3\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[3\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09104__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07729_ _03617_ _03618_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10740_ _06389_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07540__D team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10670__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10671_ net931 _04421_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12410_ net279 net2420 net488 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16776__1330 vssd1 vssd1 vccd1 vccd1 _16776__1330/HI net1330 sky130_fd_sc_hd__conb_1
X_13390_ team_02_WB.instance_to_wrap.top.a1.row1\[60\] _03226_ _03289_ _03137_ vssd1
+ vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a211o_1
XANTENNA__09812__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ net265 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] net497 vssd1
+ vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16206__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ clknet_leaf_81_wb_clk_i _01511_ _00023_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_12272_ net250 net1880 net506 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14011_ net1046 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XANTENNA__11786__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06844_ _06845_ net411 vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__mux2_1
XANTENNA__13567__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15230__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16356__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ team_02_WB.instance_to_wrap.top.pc\[18\] _06337_ vssd1 vssd1 vccd1 vccd1
+ _06781_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10703__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] net702 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\]
+ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a221o_1
X_15962_ clknet_leaf_116_wb_clk_i _02413_ _00920_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11085_ _05114_ net445 _06144_ net452 vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a22o_1
X_16732__1286 vssd1 vssd1 vccd1 vccd1 _16732__1286/HI net1286 sky130_fd_sc_hd__conb_1
X_14913_ net1149 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XANTENNA__09343__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] net853 net793 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15380__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ clknet_leaf_124_wb_clk_i _02344_ _00851_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ net1154 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XANTENNA__12410__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07504__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14775_ net1177 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11987_ net2368 net283 net533 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16514_ clknet_leaf_37_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[17\]
+ _01388_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13726_ net1018 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10938_ _04910_ net452 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__and2b_1
XANTENNA__08854__B2 team_02_WB.instance_to_wrap.ramload\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16445_ clknet_leaf_81_wb_clk_i net1696 _01319_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13657_ net1064 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
X_10869_ team_02_WB.instance_to_wrap.top.pc\[27\] _06343_ team_02_WB.instance_to_wrap.top.pc\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ _06620_ _06647_ _07235_ _06729_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__or4b_1
X_16376_ clknet_leaf_73_wb_clk_i _02807_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13588_ net1161 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XANTENNA__09803__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15327_ clknet_leaf_26_wb_clk_i _01778_ _00285_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12539_ net263 net2491 net467 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14861__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15258_ clknet_leaf_116_wb_clk_i _01709_ _00216_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11696__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14209_ net1100 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10177__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15189_ clknet_leaf_115_wb_clk_i _01640_ _00147_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09582__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 net412 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
Xfanout419 net424 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08790__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13115__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net685 net664 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08701_ _04479_ _04485_ _04491_ _04497_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09681_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] net801 net785 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__a22o_1
XANTENNA__11141__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ net910 net615 _04426_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__or3_4
XFILLER_0_20_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12320__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15873__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ net979 _04358_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net978
+ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07514_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__nor2_1
XANTENNA__13940__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _02864_ _04326_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or2_1
XANTENNA__10101__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout330_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1072_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11601__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\] net677 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15253__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09046_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] net782 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\]
+ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout797_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold440 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10168__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold451 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09573__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 team_02_WB.instance_to_wrap.ramload\[30\] vssd1 vssd1 vccd1 vccd1 net1893
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10523__B _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13106__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 _03424_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08781__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 _04403_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout942 _07365_ vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_4
X_09948_ _05595_ _05605_ _05608_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__nor4_2
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout964 net966 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 team_02_WB.instance_to_wrap.top.a1.instruction\[13\] vssd1 vssd1 vccd1
+ vccd1 net975 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 team_02_WB.instance_to_wrap.top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1
+ net986 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09325__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net998 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_2
X_09879_ _05533_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ net273 net2041 net543 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
Xhold1162 team_02_WB.instance_to_wrap.top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 net2560
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1173 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12230__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ team_02_WB.instance_to_wrap.top.pc\[5\] _05797_ vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10340__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1184 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1195 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ net261 net2391 net550 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11772_ net252 net1866 net558 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
X_14560_ net1083 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13511_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10723_ _04888_ net371 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14491_ net1060 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16230_ clknet_leaf_28_wb_clk_i _02675_ _01187_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input93_A wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ _06305_ _06240_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__nand2b_1
X_13442_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\]
+ _03303_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16161_ clknet_leaf_29_wb_clk_i net1527 _01119_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dfrtp_1
X_13373_ _03226_ _03273_ _03275_ _03272_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or4b_1
XFILLER_0_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08064__A2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net928 net590 vssd1
+ vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15112_ clknet_leaf_55_wb_clk_i _01563_ _00070_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12324_ net326 net2551 net502 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__mux2_1
XANTENNA__09775__A _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16092_ clknet_leaf_92_wb_clk_i _02538_ _01050_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15043_ net1161 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__inv_2
XANTENNA__15746__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12255_ net299 net1776 net510 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12405__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _06260_ net744 net458 team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _06829_
+ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__a221o_1
X_12186_ net285 net2123 net517 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ net400 _06420_ _06535_ _06763_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ clknet_leaf_29_wb_clk_i _02396_ _00903_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11068_ _06144_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ net462 _05545_ _05679_ net456 net740 vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12140__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15876_ clknet_leaf_19_wb_clk_i _02327_ _00834_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10331__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14827_ net1191 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
XANTENNA__15126__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14856__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ net1177 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16493__D team_02_WB.instance_to_wrap.top.aluOut\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13709_ net1130 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14689_ net1197 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11280__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15276__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ clknet_leaf_62_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[27\]
+ _01302_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire598_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16521__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16359_ clknet_leaf_101_wb_clk_i _02792_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12315__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10343__B team_02_WB.instance_to_wrap.top.DUT.read_data2\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__A2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[12\] net871 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a22o_1
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout249 _06479_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_1
X_07994_ _03841_ _03847_ _03860_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11158__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09307__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _05359_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout280_A _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12050__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09664_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] net720 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\]
+ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08615_ net973 _04373_ _04409_ _04410_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a211o_1
X_09595_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] net812 net877 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14766__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout545_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net77 net1642 net892 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15619__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11822__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ net1623 net751 net742 _04294_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout712_A _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10518__B _05521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731__1285 vssd1 vssd1 vccd1 vccd1 _16731__1285/HI net1285 sky130_fd_sc_hd__conb_1
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _05482_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\] net717 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12225__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12040_ net251 net2195 net529 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XANTENNA__09546__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\] vssd1
+ vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 net145 vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12973__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 _04424_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_2
Xfanout761 net764 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
Xfanout772 _04673_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_2
X_13991_ net1134 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
Xfanout783 _04669_ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
Xfanout794 _04661_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ clknet_leaf_10_wb_clk_i _02181_ _00688_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12942_ _02974_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10313__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15661_ clknet_leaf_24_wb_clk_i _02112_ _00619_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12873_ team_02_WB.instance_to_wrap.top.pc\[13\] _06276_ vssd1 vssd1 vccd1 vccd1
+ _02907_ sky130_fd_sc_hd__nand2_1
XANTENNA__13580__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14612_ net1193 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XANTENNA__15299__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11824_ net329 net1960 net554 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15592_ clknet_leaf_85_wb_clk_i _02043_ _00550_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16544__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14543_ net1110 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11755_ net299 net2216 net561 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XANTENNA__10709__A _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _05257_ net373 vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10092__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14474_ net1026 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11686_ net285 net1890 net568 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10428__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16213_ clknet_leaf_30_wb_clk_i _02658_ _01170_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ _03303_ _03308_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10637_ _06261_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ clknet_leaf_38_wb_clk_i net1546 _01102_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10568_ net929 _04628_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and2b_2
XFILLER_0_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13356_ team_02_WB.instance_to_wrap.top.a1.row2\[42\] _03230_ _03239_ team_02_WB.instance_to_wrap.top.a1.row1\[122\]
+ _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ net258 net1850 net501 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__mux2_1
X_16075_ clknet_leaf_22_wb_clk_i _02526_ _01033_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13287_ _03179_ _03185_ _03196_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__o211ai_1
XANTENNA__10444__A _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ _05402_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09537__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15026_ net1154 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ net247 net1925 net509 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08745__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net238 net2338 net516 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap608_A _05480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16488__D team_02_WB.instance_to_wrap.top.aluOut\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16074__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 wb_rst_i vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16755__1309 vssd1 vssd1 vccd1 vccd1 _16755__1309/HI net1309 sky130_fd_sc_hd__conb_1
X_15928_ clknet_leaf_121_wb_clk_i _02379_ _00886_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10304__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09170__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ clknet_leaf_126_wb_clk_i _02310_ _00817_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12057__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ net1669 net935 net918 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1
+ vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
X_09380_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\] net821 net761 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08331_ _04205_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07484__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08262_ _04123_ _04136_ _04126_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08193_ _04045_ _04057_ net224 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__and3_1
XANTENNA__13021__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12045__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07977_ _03858_ _03859_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1
+ vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout662_A _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11185__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09716_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[14\] net813 net810 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16567__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ _05296_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] net663 net650 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12599__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ net96 net1611 net891 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XANTENNA__15591__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07475__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11540_ net356 net2256 net585 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XANTENNA__10074__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11271__B2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire425 _07280_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_1
X_11471_ net913 _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12744__A _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13026__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ team_02_WB.START_ADDR_VAL_REG\[18\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net201 sky130_fd_sc_hd__a21o_1
XANTENNA__11023__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ net580 net373 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nor2_1
XANTENNA__09767__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ net1116 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _03134_
+ sky130_fd_sc_hd__nand3_1
X_10353_ _05884_ _06003_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and2b_1
XANTENNA__07557__B team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09519__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ team_02_WB.instance_to_wrap.top.pc\[10\] _05593_ vssd1 vssd1 vccd1 vccd1
+ _03085_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input56_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10284_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\] net869 net781 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a221o_1
XANTENNA__12523__A1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08727__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net301 net2480 net469 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
XANTENNA__13575__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout580 _04624_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
Xfanout591 _06221_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16762_ net1316 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
X_13974_ net1109 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XANTENNA__09152__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15713_ clknet_leaf_2_wb_clk_i _02164_ _00671_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ _02958_ _02898_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__nand2b_1
X_16693_ net1247 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15934__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15644_ clknet_leaf_63_wb_clk_i _02095_ _00602_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ team_02_WB.instance_to_wrap.top.pc\[23\] _06246_ vssd1 vssd1 vccd1 vccd1
+ _02890_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net260 net2384 net555 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
X_15575_ clknet_leaf_118_wb_clk_i _02026_ _00533_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12787_ _05889_ _05929_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14526_ net1022 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XANTENNA__11262__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ net249 net2672 net562 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10158__B team_02_WB.instance_to_wrap.top.DUT.read_data2\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14457_ net1059 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
X_11669_ net240 net2275 net570 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13003__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15030__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ net1473 _04236_ net828 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09758__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ net1052 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ clknet_leaf_65_wb_clk_i _02573_ _01085_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13339_ net985 _03212_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nand2_1
X_16058_ clknet_leaf_123_wb_clk_i _02509_ _01016_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08718__B1 _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ net1163 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__inv_2
X_07900_ _03743_ _03755_ _03784_ _03742_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a22o_2
XFILLER_0_62_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ net959 _04315_ _04328_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] vssd1
+ vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a22o_1
XANTENNA__15464__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ _03682_ _03719_ _03721_ _03710_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16730__1284 vssd1 vssd1 vccd1 vccd1 _16730__1284/HI net1284 sky130_fd_sc_hd__conb_1
X_07762_ _03613_ _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09501_ _05158_ _05159_ _05171_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or4_4
XFILLER_0_116_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07693_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03541_ net362 vssd1 vssd1
+ vccd1 vccd1 _03584_ sky130_fd_sc_hd__or3b_1
XFILLER_0_91_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09432_ _05100_ _05102_ _05104_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09363_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\] net698 _05038_ vssd1
+ vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10056__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _04170_ _04171_ _04175_ _04182_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or4b_1
X_09294_ _04962_ _04971_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__nor2_8
XANTENNA_10 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ _04124_ _04125_ _04121_ _04122_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11879__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08176_ net2640 net936 net920 net224 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09749__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11556__A2 _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10084__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[8] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[17] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout877_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[8] sky130_fd_sc_hd__buf_2
XANTENNA__12503__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XANTENNA__09382__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15957__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09134__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10971_ _06239_ _06240_ _06305_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _05936_ _05975_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10295__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ net1046 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12641_ _06145_ _06186_ _07267_ _07268_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__or4_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10047__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15360_ clknet_leaf_9_wb_clk_i _01811_ _00318_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12572_ net263 net1785 net474 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__mux2_1
XANTENNA__09988__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08952__A team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ net1136 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15337__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__B2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ _05836_ net374 _06109_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__a21oi_1
X_15291_ clknet_leaf_105_wb_clk_i _01742_ _00249_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242_ net1091 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11454_ net426 _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16754__1308 vssd1 vssd1 vccd1 vccd1 _16754__1308/HI net1308 sky130_fd_sc_hd__conb_1
XFILLER_0_22_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10706__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10405_ _05175_ net367 vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__nand2_1
XANTENNA__12624__D _06629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ team_02_WB.instance_to_wrap.top.pc\[10\] net907 _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a221o_1
X_14173_ net1031 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ net1596 _03126_ _03127_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a21bo_1
X_10336_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\] net807 net799 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a22o_1
X_10267_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] net685 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13055_ _07395_ _07396_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__nor2_1
XANTENNA__12413__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ net248 net2641 net470 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__mux2_1
XANTENNA__09373__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] net872 net804 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\]
+ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11180__B1 team_02_WB.instance_to_wrap.top.aluOut\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16814_ net1368 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16745_ net1299 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
XFILLER_0_89_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13957_ net1074 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
X_12908_ _02939_ _02941_ _02914_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10286__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16676_ net1230 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ net1070 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_128_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15627_ clknet_leaf_21_wb_clk_i _02078_ _00585_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12839_ _04723_ _06223_ _02872_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14864__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09979__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ clknet_leaf_12_wb_clk_i _02009_ _00516_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11699__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ net1132 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15489_ clknet_leaf_129_wb_clk_i _01940_ _00447_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08030_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__inv_2
Xinput30 wbm_dat_i[30] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_126_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput52 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12735__A1 _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold803 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold814 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
Xinput85 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xhold825 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xinput96 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_1
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold847 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold858 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold869 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] net803 net787 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\]
+ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08932_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] net653 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12323__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09364__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ net1600 _04559_ net825 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
XANTENNA__10351__B _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ net341 _03679_ _03654_ _03658_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08794_ net171 net953 net904 net1494 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09116__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ _03621_ _03632_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout458_A _06326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _03535_ _03564_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] net685 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16605__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13215__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _05016_ _05018_ _05020_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09277_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] net706 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\]
+ _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ _04064_ _04070_ _04081_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08159_ _04020_ _04023_ _04032_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10201__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ net405 _06575_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12741__B team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\] net835 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ _05779_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12233__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _05705_ _05707_ _05709_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14860_ net1174 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XANTENNA__09107__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ net1144 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XANTENNA_input19_A wbm_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14791_ net1173 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16530_ clknet_leaf_74_wb_clk_i _02828_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13742_ net1063 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XANTENNA__10268__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ net391 _06454_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16461_ clknet_leaf_65_wb_clk_i net1544 _01335_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13673_ net1028 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
X_10885_ _06528_ _06529_ net403 vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15412_ clknet_leaf_51_wb_clk_i _01863_ _00370_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ _06532_ _06577_ _06597_ _06629_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__or4_1
X_16392_ clknet_leaf_77_wb_clk_i _02823_ _01266_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15343_ clknet_leaf_32_wb_clk_i _01794_ _00301_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12555_ net326 net2419 net465 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__mux2_1
XANTENNA__12408__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10976__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11506_ net422 _06733_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15274_ clknet_leaf_43_wb_clk_i _01725_ _00232_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12486_ net301 net1816 net482 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ net1031 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
X_11437_ net416 _07041_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09594__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ net1005 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ _06385_ _06390_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13107_ net231 _03112_ _03113_ _07419_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12143__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] net703 net696 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a221o_1
X_14087_ net1153 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XANTENNA__10452__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11299_ _06088_ _06090_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__nand2_1
X_13038_ net231 _03055_ net228 _06836_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09018__A _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11982__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14859__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13763__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1169 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_4
Xfanout1172 net1185 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_4
Xfanout1183 net1184 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16496__D team_02_WB.instance_to_wrap.top.aluOut\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14989_ net1173 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
XANTENNA__15502__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ _03419_ net936 vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16728_ net1282 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07461_ team_02_WB.instance_to_wrap.top.pc\[20\] vssd1 vssd1 vccd1 vccd1 _03402_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ net1393 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_130_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] net683 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\]
+ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09688__A _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] net818 net774 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\]
+ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a221o_1
XANTENNA__12956__B2 _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12318__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09062_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] net700 net641 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10346__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08013_ _03871_ net241 _03898_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a22oi_4
XANTENNA__16008__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold600 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold622 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold633 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold655 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold666 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold677 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\] net670 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a22o_1
XANTENNA__12053__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16158__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09337__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__inv_2
X_09895_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\] net779 _05558_ vssd1
+ vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout575_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 team_02_WB.START_ADDR_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11892__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1311 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ net10 net948 net922 net1786 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__o22a_1
Xhold1333 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1344 team_02_WB.instance_to_wrap.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net2742
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15182__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ net1590 net956 net927 _04545_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
X_16753__1307 vssd1 vssd1 vccd1 vccd1 _16753__1307/HI net1307 sky130_fd_sc_hd__conb_1
XFILLER_0_79_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07659_ _03509_ _03537_ _03522_ _03517_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_32_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] _06321_ _04583_ vssd1 vssd1
+ vccd1 vccd1 _06322_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ _04998_ _05003_ _05004_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or4_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12228__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ net260 net1992 net496 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12271_ net246 net2396 net506 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux2_1
XANTENNA__12752__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ net1053 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11222_ _06622_ _06624_ net404 vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09040__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ net305 net1965 net585 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09328__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\] net657 net637 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a22o_1
X_11084_ net435 _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__nor2_1
X_15961_ clknet_leaf_108_wb_clk_i _02412_ _00919_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14912_ net1159 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XANTENNA__13583__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\] net878 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a221o_1
X_15892_ clknet_leaf_51_wb_clk_i _02343_ _00850_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ net1161 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ net1178 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
X_11986_ net2142 net267 net532 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09500__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16513_ clknet_leaf_0_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[16\]
+ _01387_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13725_ net1105 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XANTENNA__10110__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10937_ net448 _06412_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08854__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10110__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16444_ clknet_leaf_81_wb_clk_i net1467 _01318_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13656_ net1056 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ net440 _06481_ _06514_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[28\]
+ sky130_fd_sc_hd__o21bai_4
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ _06588_ _07234_ _06676_ _06701_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__or4b_1
XFILLER_0_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16375_ clknet_leaf_73_wb_clk_i _02806_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12138__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ net1161 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10799_ net384 _06442_ _06446_ _06447_ net393 vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__o221a_1
XFILLER_0_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ clknet_leaf_6_wb_clk_i _01777_ _00284_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12538_ net260 net2254 net467 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11977__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15257_ clknet_leaf_106_wb_clk_i _01708_ _00215_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12469_ net246 net1904 net481 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14208_ net1082 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_15188_ clknet_leaf_51_wb_clk_i _01639_ _00146_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09031__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ net1048 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout409 net412 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] net622 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09680_ _05342_ _05344_ _05346_ _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08631_ net910 net615 _04426_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nor3_4
XFILLER_0_59_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11429__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04358_ vssd1 vssd1 vccd1
+ vccd1 _04359_ sky130_fd_sc_hd__nand2_1
XANTENNA__11429__B2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09098__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07513_ net2432 net117 _00011_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ team_02_WB.instance_to_wrap.top.a1.row1\[63\] _04325_ _04329_ vssd1 vssd1
+ vccd1 vccd1 _02684_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08845__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12048__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[28\] net669 net641 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09270__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11887__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[30\] net813 net845 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold430 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09022__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold441 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] vssd1
+ vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold485 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold496 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout910 _04384_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_4
XFILLER_0_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_2
XANTENNA__08781__B2 _04547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09947_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\] net791 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\]
+ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a221o_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
Xfanout954 _04340_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 team_02_WB.instance_to_wrap.top.a1.instruction\[12\] vssd1 vssd1 vccd1
+ vccd1 net976 sky130_fd_sc_hd__buf_2
XANTENNA__12511__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _05535_ _05537_ _05539_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1
+ net987 sky130_fd_sc_hd__clkbuf_2
Xfanout998 net61 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_2
Xhold1130 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08829_ net28 net947 net921 net1707 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__o22a_1
Xhold1152 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net255 net1948 net550 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11771_ net247 net1869 net558 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08836__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__A _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13510_ team_02_WB.instance_to_wrap.top.pad.button_control.debounce team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10722_ _04932_ net373 vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_1
X_14490_ net1058 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13441_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] _03303_ net1676 vssd1 vssd1
+ vccd1 vccd1 _03319_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10653_ team_02_WB.instance_to_wrap.top.pc\[24\] _06242_ _06304_ vssd1 vssd1 vccd1
+ vccd1 _06305_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16160_ clknet_leaf_37_wb_clk_i net1482 _01118_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input86_A wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13372_ _03397_ team_02_WB.instance_to_wrap.top.lcd.nextState\[4\] _03212_ _03274_
+ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10584_ team_02_WB.instance_to_wrap.top.pc\[26\] _06234_ vssd1 vssd1 vccd1 vccd1
+ _06236_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09261__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11797__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ clknet_leaf_13_wb_clk_i _01562_ _00069_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net313 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\] net502 vssd1
+ vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XANTENNA__13578__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16091_ clknet_leaf_93_wb_clk_i _02537_ _01049_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09549__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ net1158 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__inv_2
X_12254_ net291 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\] net508 vssd1
+ vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__mux2_1
X_11205_ net914 _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ net269 net1857 net516 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ net416 _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12421__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _05154_ _06033_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__or2_1
X_15944_ clknet_leaf_56_wb_clk_i _02395_ _00902_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07515__S _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] net615 _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a22o_2
X_15875_ clknet_leaf_43_wb_clk_i _02326_ _00833_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14826_ net1192 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
XANTENNA__09015__B _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14757_ net1181 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XANTENNA__08827__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11969_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04576_ _07187_ _07204_
+ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10095__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15033__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ net1018 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
X_14688_ net1197 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ net1135 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
X_16427_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[26\]
+ _01301_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09788__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_102_wb_clk_i _02791_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15309_ clknet_leaf_22_wb_clk_i _01760_ _00267_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16289_ clknet_leaf_94_wb_clk_i _02722_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfxtp_1
X_16752__1306 vssd1 vssd1 vccd1 vccd1 _16752__1306/HI net1306 sky130_fd_sc_hd__conb_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639__1210 vssd1 vssd1 vccd1 vccd1 _16639__1210/HI net1210 sky130_fd_sc_hd__conb_1
XANTENNA__13336__B2 team_02_WB.instance_to_wrap.top.a1.row2\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09801_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] net821 net819 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08763__B2 _04538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09960__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 _07336_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_4
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_07993_ _03841_ _03842_ _03846_ _03860_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__and4_1
XANTENNA__10570__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _05378_ _05397_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__nor2_1
XANTENNA__12331__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09712__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\] net704 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout273_A _06674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ net976 _04379_ _04406_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\] net784 net756 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ net78 net1631 net892 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08818__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11471__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15220__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16346__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08476_ net1588 net751 net742 _04291_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09491__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout705_A _04461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09779__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15370__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16496__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12506__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _04705_ _04707_ _04709_ _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__or4_4
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 team_02_WB.instance_to_wrap.top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1 net1658
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_02_WB.instance_to_wrap.top.a1.row2\[0\] vssd1 vssd1 vccd1 vccd1 net1669
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_02_WB.instance_to_wrap.top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 net1680
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold293 _02804_ vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_2
Xfanout751 _04323_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
Xfanout762 net764 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XANTENNA__12241__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout773 _04671_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14022__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ net1139 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
Xfanout784 _04669_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_2
Xfanout795 _04661_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09703__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ team_02_WB.instance_to_wrap.top.pc\[31\] _06222_ vssd1 vssd1 vccd1 vccd1
+ _02975_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15660_ clknet_leaf_52_wb_clk_i _02111_ _00618_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ team_02_WB.instance_to_wrap.top.pc\[15\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _02906_ sky130_fd_sc_hd__xnor2_1
X_14611_ net1196 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11823_ net313 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net554 vssd1
+ vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
X_15591_ clknet_leaf_14_wb_clk_i _02042_ _00549_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10077__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ net1116 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ net293 net2380 net560 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10705_ _06352_ _06355_ net364 vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ net1025 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
X_11685_ net270 net2117 net568 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ clknet_leaf_28_wb_clk_i _02657_ _01169_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13424_ net994 _03303_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__and3_1
X_10636_ team_02_WB.instance_to_wrap.top.pc\[17\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _06288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16143_ clknet_leaf_128_wb_clk_i net1577 _01101_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13355_ team_02_WB.instance_to_wrap.top.a1.row1\[114\] _03219_ _03234_ team_02_WB.instance_to_wrap.top.a1.row2\[18\]
+ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a22o_1
XANTENNA__10725__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12416__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ net441 _06054_ net429 _06219_ _06138_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[31\]
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11320__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ net256 net2590 net500 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__mux2_1
X_16074_ clknet_leaf_45_wb_clk_i _02525_ _01032_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13286_ _03178_ _03191_ _03184_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10444__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498_ _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__nor2_2
XFILLER_0_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15025_ net1154 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12237_ net242 net2442 net508 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10001__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__B2 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12168_ _04576_ _04579_ _07190_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12767__A_N _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16219__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ net912 _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__nor2_1
XANTENNA__12151__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net352 net2019 net524 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput6 wbm_ack_i vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
X_15927_ clknet_leaf_118_wb_clk_i _02378_ _00885_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11990__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ clknet_leaf_25_wb_clk_i _02309_ _00816_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14809_ net1203 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15789_ clknet_leaf_43_wb_clk_i _02240_ _00747_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10068__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ _04186_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08261_ _04136_ _04138_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08192_ _04057_ net224 _04075_ _04074_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09225__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12326__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09933__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _03830_ _03860_ _03864_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_96_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09715_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\] net858 net850 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09646_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[16\] net592 vssd1
+ vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09577_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\] net735 net723 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a22o_1
XANTENNA__15736__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08528_ _04345_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09464__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11271__A2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ team_02_WB.instance_to_wrap.top.a1.data\[2\] net916 vssd1 vssd1 vccd1 vccd1
+ _04314_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15886__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11470_ team_02_WB.instance_to_wrap.top.pc\[6\] _06329_ vssd1 vssd1 vccd1 vccd1 _07072_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09216__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10421_ _04804_ net368 _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12236__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13140_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ net398 _05883_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__nand2_1
XANTENNA__07557__C team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15116__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13071_ team_02_WB.instance_to_wrap.top.pc\[11\] net945 net941 _03084_ vssd1 vssd1
+ vccd1 vccd1 _01509_ sky130_fd_sc_hd__a22o_1
X_10283_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[1\] net861 net805 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__a22o_1
XANTENNA__12760__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09924__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ net291 net2362 net468 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XANTENNA_input49_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A0 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout570 _07193_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout592 _04631_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
X_13973_ net1120 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
X_16761_ net1315 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08509__A_N net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10298__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ team_02_WB.instance_to_wrap.top.pc\[19\] _06257_ _02957_ vssd1 vssd1 vccd1
+ vccd1 _02958_ sky130_fd_sc_hd__a21o_1
X_15712_ clknet_leaf_10_wb_clk_i _02163_ _00670_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_16692_ net1246 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12855_ team_02_WB.instance_to_wrap.top.pc\[23\] _06246_ vssd1 vssd1 vccd1 vccd1
+ _02889_ sky130_fd_sc_hd__and2_1
X_15643_ clknet_leaf_118_wb_clk_i _02094_ _00601_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_16751__1305 vssd1 vssd1 vccd1 vccd1 _16751__1305/HI net1305 sky130_fd_sc_hd__conb_1
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11806_ net254 net1821 net553 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15574_ clknet_leaf_109_wb_clk_i _02025_ _00532_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ _05887_ _05888_ _05929_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09455__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14525_ net1031 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
X_11737_ net244 net2525 net562 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08663__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14456_ net1056 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
X_11668_ _04428_ _04579_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__or3_4
XFILLER_0_25_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ net1476 _04245_ net828 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
X_10619_ net750 _05886_ _06270_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__o21a_2
XANTENNA__10455__A _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12146__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net1128 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
X_11599_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] _04428_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__or3b_2
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16126_ clknet_leaf_64_wb_clk_i _02572_ _01084_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10222__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ net2322 net895 _03243_ net993 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o211a_1
XANTENNA__16041__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13766__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ clknet_leaf_107_wb_clk_i _02508_ _01015_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13269_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[1\] team_02_WB.instance_to_wrap.top.pad.keyCode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__or4b_2
XFILLER_0_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08718__A1 _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ net1163 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16499__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07830_ _03717_ _03718_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07761_ _03612_ net350 vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15759__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] net727 net714 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\]
+ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a221o_1
XANTENNA__10289__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07692_ _03407_ net362 _03541_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09694__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] net865 net814 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09362_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\] net714 net642 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09446__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ _04172_ _04179_ _04181_ _04175_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09293_ _04964_ _04966_ _04968_ _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__or4_2
XANTENNA__08654__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A _07186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _04124_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08534__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ _04039_ _04059_ _04035_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12056__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1145_A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10764__A1 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11895__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[28] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08709__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[18] sky130_fd_sc_hd__buf_2
XANTENNA__08709__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09906__B1 _05568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[9] sky130_fd_sc_hd__buf_2
X_16655__1389 vssd1 vssd1 vccd1 vccd1 net1389 _16655__1389/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout772_A _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__11196__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07959_ _03842_ _03845_ _03846_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ _06609_ _06610_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[25\]
+ sky130_fd_sc_hd__or2_2
XANTENNA__09685__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12739__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] net869 net789 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12640_ _04703_ _06142_ _06143_ net452 vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__or4b_1
XFILLER_0_116_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input103_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ net258 net1809 net474 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__mux2_1
XANTENNA__08951__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__B team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14310_ net1092 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11522_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] net887 net907 team_02_WB.instance_to_wrap.top.pc\[3\]
+ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15290_ clknet_leaf_123_wb_clk_i _01741_ _00248_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14241_ net1100 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
X_11453_ _05749_ _06164_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10404_ _04601_ _06055_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or2_1
X_14172_ net1098 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11384_ net913 _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _03126_ net990 _04274_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__or3b_1
X_10335_ _05982_ _05984_ _05986_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07584__A team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13154__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13054_ net230 _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__nand2_1
X_10266_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\] net672 net644 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10722__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ net243 net1932 net470 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10197_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\] net852 net844 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a22o_1
XANTENNA__11180__A1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16813_ net1367 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11834__A team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16744_ net1298 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13956_ net1141 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__09676__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12907_ _02914_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13887_ net1118 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16675_ team_02_WB.instance_to_wrap.top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 net107
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15626_ clknet_leaf_44_wb_clk_i _02077_ _00584_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12838_ _07368_ _02871_ _07367_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09428__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15557_ clknet_leaf_126_wb_clk_i _02008_ _00515_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12769_ _05378_ _06268_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14508_ net1004 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
X_15488_ clknet_leaf_11_wb_clk_i _01939_ _00446_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 wbm_dat_i[21] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput31 wbm_dat_i[31] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1152 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_1
Xinput53 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09974__A _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15431__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xinput75 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput86 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold815 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
Xhold837 team_02_WB.instance_to_wrap.top.pc\[15\] vssd1 vssd1 vccd1 vccd1 net2235
+ sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ clknet_leaf_64_wb_clk_i _02555_ _01067_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold848 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] net859 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10913__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold859 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] net706 net674 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\]
+ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15581__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net959 _04290_ _04302_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a32o_1
X_07813_ net341 _03679_ _03654_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__a21oi_1
X_08793_ net172 net953 net904 net1481 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07744_ _03621_ _03632_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08529__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07675_ _03562_ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and2_1
XANTENNA__12671__A1 _06963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout353_A _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1095_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] net736 net676 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] net792 net840 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[23\]
+ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout520_A _07212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12974__A2 _07336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\] net713 net674 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08227_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04028_ _04071_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__or4b_1
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_107_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09052__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ _04041_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12514__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15924__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _03950_ net225 _03939_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a21oi_1
X_16750__1304 vssd1 vssd1 vccd1 vccd1 _16750__1304/HI net1304 sky130_fd_sc_hd__conb_1
XFILLER_0_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] net871 net851 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a22o_1
X_10051_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] net686 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ _05710_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a221o_1
XANTENNA__13151__A2 _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ net1080 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
X_14790_ net1177 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ net1134 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10953_ _06451_ _06453_ net390 vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16460_ clknet_leaf_64_wb_clk_i net1659 _01334_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13672_ net1096 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
X_10884_ net390 _06115_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08963__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15411_ clknet_leaf_124_wb_clk_i _01862_ _00369_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12623_ _06219_ _06431_ _07250_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16391_ clknet_leaf_77_wb_clk_i _02822_ _01265_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11217__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15342_ clknet_leaf_41_wb_clk_i _01793_ _00300_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12554_ net311 net2639 net464 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__mux2_1
XANTENNA__15454__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09291__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10976__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10976__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06008_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15273_ clknet_leaf_29_wb_clk_i _01724_ _00231_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12485_ net293 net2120 net480 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ net1018 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11436_ net393 _06874_ _07039_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__o22a_1
XANTENNA__09043__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11925__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13390__A2 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ net1014 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XANTENNA__12424__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ _05572_ _06018_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _07409_ _07416_ _07418_ net890 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__o31ai_1
X_10318_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\] net706 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a22o_1
X_14086_ net1140 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
X_11298_ net400 _06711_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__nand2_1
XANTENNA__10452__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13037_ _07390_ _07441_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10249_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] net857 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a22o_1
XANTENNA__09018__B _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_2
XANTENNA__09897__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1151 net1160 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1162 net1165 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_4
Xfanout1173 net1185 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1204 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_2
X_14988_ net1191 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16727_ net1281 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__11283__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ net1128 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
X_07460_ team_02_WB.instance_to_wrap.top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16658_ net1392 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_53_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15609_ clknet_leaf_117_wb_clk_i _02060_ _00567_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10908__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16589_ clknet_leaf_58_wb_clk_i net1405 _01462_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654__1388 vssd1 vssd1 vccd1 vccd1 net1388 _16654__1388/LO sky130_fd_sc_hd__conb_1
X_09130_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\] net843 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _04742_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08012_ _03827_ _03870_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold601 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold612 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold623 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold634 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold656 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 team_02_WB.instance_to_wrap.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2065
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09209__A _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] net722 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a221o_1
Xhold678 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ net976 _04407_ _04409_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09894_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\] net880 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1010_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1301 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ net11 net948 net922 net2239 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__o22a_1
Xhold1312 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1323 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1334 team_02_WB.instance_to_wrap.top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1
+ net2732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1345 team_02_WB.instance_to_wrap.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net2743
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout568_A _07193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08776_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[4\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[4\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_2
XFILLER_0_58_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07727_ _03589_ _03609_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14785__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout735_A _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07658_ _03509_ _03537_ _03517_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15477__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ _03447_ _03450_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\] net651 net627 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ _04999_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09812__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\] net820 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[25\]
+ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12270_ net244 net2394 net506 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08722__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11221_ net404 _06625_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12244__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11152_ net460 team_02_WB.instance_to_wrap.top.aluOut\[19\] _06777_ _06779_ vssd1
+ vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__o22a_2
XFILLER_0_43_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10103_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] net726 net682 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15960_ clknet_leaf_121_wb_clk_i _02411_ _00918_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11083_ net416 _06715_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__or2_1
XANTENNA__08958__A team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A wbm_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ net1162 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
X_10034_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] net849 net777 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a22o_1
X_15891_ clknet_leaf_124_wb_clk_i _02342_ _00849_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11384__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1161 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08839__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11985_ net2727 net323 net532 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
X_14773_ net1177 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16512_ clknet_leaf_7_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[15\]
+ _01386_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10936_ _06578_ net413 net436 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__and3b_1
X_13724_ net1097 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16443_ clknet_leaf_91_wb_clk_i net1574 _01317_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13655_ net1107 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XANTENNA__12419__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ net428 _06482_ _06500_ net439 _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ _06755_ _06787_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16374_ clknet_leaf_73_wb_clk_i _02805_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13586_ net1154 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ net378 _06074_ net388 vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09803__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12537_ net254 net2599 net466 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15325_ clknet_leaf_111_wb_clk_i _01776_ _00283_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12468_ net244 net2468 net481 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
X_15256_ clknet_leaf_122_wb_clk_i _01707_ _00214_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14207_ net1121 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
X_11419_ _04625_ net407 _07024_ _07025_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__a31o_1
X_15187_ clknet_leaf_126_wb_clk_i _01638_ _00145_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12154__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ net236 net2018 net494 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10177__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14138_ net1053 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11993__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13115__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ net1117 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
X_16821__1375 vssd1 vssd1 vccd1 vccd1 _16821__1375/HI net1375 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _04367_ _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__or2_2
XFILLER_0_94_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ team_02_WB.instance_to_wrap.top.a1.instruction\[2\] team_02_WB.instance_to_wrap.top.a1.instruction\[1\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[0\] vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07512_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__and2b_1
XFILLER_0_136_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07502__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ _04327_ _04280_ _04279_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10101__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_112_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12329__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13051__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] net665 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12853__A team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1058_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\] net767 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold420 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13354__A2 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold431 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10168__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold442 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold464 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold475 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xfanout922 _04556_ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[9\] net876 net842 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout944 _07363_ vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_2
Xfanout955 net958 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_2
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_2
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
Xhold1120 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout852_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[10\] net738 net705 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\]
+ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a221o_1
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10876__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout999 net1015 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09730__A1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1142 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08828_ net30 net949 net923 net1893 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
Xhold1153 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10340__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ net1585 net957 net925 _04536_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
Xhold1197 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ net244 net2135 net558 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA__09494__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10721_ net378 _06370_ _06371_ _06369_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12239__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13440_ net1678 _03303_ _03318_ net1176 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a211oi_1
X_10652_ _06243_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__and2_1
XANTENNA__09246__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13371_ _03215_ _03231_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12763__A _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ net307 net2232 net503 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15110_ clknet_leaf_11_wb_clk_i _01561_ _00068_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16090_ clknet_leaf_80_wb_clk_i _02536_ _01048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input79_A wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15041_ net1156 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12253_ net285 net2690 net508 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XANTENNA__16618__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__A2 _05797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11204_ _06337_ _06827_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ net323 net2625 net516 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11135_ net400 _06539_ _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11108__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15943_ clknet_leaf_14_wb_clk_i _02394_ _00901_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11066_ net281 net2213 net584 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _05677_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10867__B1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15874_ clknet_leaf_47_wb_clk_i _02325_ _00832_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10331__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14825_ net1192 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
XANTENNA__15792__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09485__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ net1179 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
X_11968_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ _04429_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11292__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ net1026 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XANTENNA__12149__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ _04913_ _06206_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__xnor2_1
X_14687_ net1196 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10458__A _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ net358 net1799 net544 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ clknet_leaf_62_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[25\]
+ _01300_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16148__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09237__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13638_ net1092 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11988__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16357_ clknet_leaf_101_wb_clk_i _02790_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ net1171 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11595__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15308_ clknet_leaf_23_wb_clk_i _01759_ _00266_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16288_ clknet_leaf_96_wb_clk_i _02721_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15172__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15239_ clknet_leaf_14_wb_clk_i _01690_ _00197_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08763__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\] net855 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07992_ _03863_ _03872_ _03873_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o31a_1
Xfanout229 net232 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10570__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__A_N _05503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\] net688 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08613_ net976 _04364_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__nor2_1
X_09593_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] net791 net840 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\]
+ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_A _06618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08544_ net79 net1665 net891 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09476__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08475_ net1627 net752 _04324_ _04288_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a22o_1
XANTENNA__12059__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1175_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11898__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold1283_A team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09027_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\] net658 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\]
+ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15665__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold250 team_02_WB.instance_to_wrap.top.a1.instruction\[1\] vssd1 vssd1 vccd1 vccd1
+ net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 team_02_WB.instance_to_wrap.top.pc\[27\] vssd1 vssd1 vccd1 vccd1 net1659
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 team_02_WB.START_ADDR_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 net130 vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_02_WB.instance_to_wrap.ramload\[24\] vssd1 vssd1 vccd1 vccd1 net1692
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A1 _04627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_8
Xfanout741 _04423_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ net456 _04509_ _05546_ net463 net740 vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a221o_1
Xfanout752 _04323_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_2
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_6
Xfanout774 _04671_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_4
Xfanout785 net788 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_8
Xfanout796 _04661_ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12940_ _02876_ _02973_ _02877_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10313__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12871_ team_02_WB.instance_to_wrap.top.pc\[16\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _02905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14610_ net1194 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
X_11822_ net307 net1876 net555 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__mux2_1
XANTENNA__09467__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15590_ clknet_leaf_13_wb_clk_i _02041_ _00548_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14541_ net1131 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11753_ net284 net1889 net562 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10704_ _06353_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09219__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11684_ net325 net2375 net568 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__mux2_1
X_14472_ net1090 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ clknet_leaf_30_wb_clk_i _02656_ _01168_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ _06284_ _06286_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nor2_1
X_16820__1374 vssd1 vssd1 vccd1 vccd1 _16820__1374/HI net1374 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16440__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ clknet_leaf_128_wb_clk_i net1491 _01100_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13354_ team_02_WB.instance_to_wrap.top.a1.row1\[58\] _03226_ _03235_ team_02_WB.instance_to_wrap.top.a1.row2\[2\]
+ _03255_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ _06217_ _06218_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__nor2_1
XANTENNA__10725__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ net250 net2585 net500 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13285_ _03185_ _03188_ _03195_ _03174_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__o211a_1
X_16073_ clknet_leaf_29_wb_clk_i _02524_ _01031_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11329__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10497_ _05484_ _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or2_1
X_12236_ net237 net2418 net508 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__mux2_1
X_15024_ net1154 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12432__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ net234 net1802 net523 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10741__A _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11118_ _06339_ _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12098_ net355 net2199 net527 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11049_ net414 _06683_ _06411_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__a21o_1
X_15926_ clknet_leaf_111_wb_clk_i _02377_ _00884_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 wbm_dat_i[0] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10304__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09170__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ clknet_leaf_19_wb_clk_i _02308_ _00815_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14808_ net1183 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XANTENNA__09458__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15788_ clknet_leaf_52_wb_clk_i _02239_ _00746_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14739_ net1200 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _04135_ _04136_ _04129_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16409_ clknet_leaf_69_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[8\]
+ _01283_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] sky130_fd_sc_hd__dfrtp_4
X_08191_ _04019_ _04054_ _04056_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15688__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12342__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07975_ _03858_ _03859_ _03831_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_103_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout383_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net798 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a22o_1
XANTENNA__09161__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ _05307_ _05311_ _05313_ _05314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[16\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_74_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout550_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout648_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ _05240_ _05242_ _05244_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__or4_4
XANTENNA__09449__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ _03412_ net933 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__nor2_2
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14793__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _04313_ net1743 net827 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08389_ _04257_ _04258_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__a21o_1
XANTENNA__12517__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _04764_ net368 vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09621__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10351_ net398 _05883_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ net230 _03080_ _03083_ net890 _03081_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a221o_1
XANTENNA__08730__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10282_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\] net761 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12021_ net283 net2533 net470 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12252__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout560 net563 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_8
Xfanout571 _07193_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16760_ net1314 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
Xfanout582 _04580_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_6
X_13972_ net1036 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
Xfanout593 _04631_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09152__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15711_ clknet_leaf_27_wb_clk_i _02162_ _00669_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12923_ _02899_ _02956_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16691_ net1245 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15642_ clknet_leaf_122_wb_clk_i _02093_ _00600_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12854_ team_02_WB.instance_to_wrap.top.pc\[24\] _04629_ vssd1 vssd1 vccd1 vccd1
+ _02888_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ net251 net2512 net553 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15573_ clknet_leaf_116_wb_clk_i _02024_ _00531_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12785_ _05843_ _05883_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14524_ net1098 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
X_11736_ net238 net2691 net562 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ net1111 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11667_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ _04428_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1
+ _07192_ sky130_fd_sc_hd__or4b_1
XANTENNA__12427__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13406_ net1507 _04253_ net828 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
X_10618_ net931 _04507_ _06220_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11598_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] _04429_ vssd1 vssd1 vccd1
+ vccd1 _07187_ sky130_fd_sc_hd__and2_1
XANTENNA__09612__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14386_ net1085 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XANTENNA__08415__B2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10455__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16125_ clknet_leaf_64_wb_clk_i _02571_ _01083_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13337_ team_02_WB.instance_to_wrap.top.a1.row2\[40\] _03230_ _03236_ _03242_ _03229_
+ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__a2111o_1
X_10549_ _04993_ _06201_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__and2b_1
XANTENNA__15980__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ clknet_leaf_121_wb_clk_i _02507_ _01014_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13268_ _03178_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__nor2_1
X_15007_ net1191 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12162__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ net268 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[15\] net512 vssd1
+ vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13199_ team_02_WB.START_ADDR_VAL_REG\[7\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net221 sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15210__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09391__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14878__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ _03612_ _03613_ net350 vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_97_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09679__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ clknet_leaf_128_wb_clk_i _02360_ _00867_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_07691_ _03407_ net362 vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09430_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net869 net861 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09361_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\] net690 net682 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\]
+ _05036_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08312_ _04172_ _04182_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\] net677 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\]
+ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08243_ _04068_ _04100_ _04119_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12337__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _04045_ _04049_ _04057_ _04042_ _04041_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09603__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[29] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 wbm_cyc_o sky130_fd_sc_hd__buf_2
XANTENNA__09906__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__12072__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__A _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 wbm_sel_o[0] sky130_fd_sc_hd__buf_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__09382__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15703__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07958_ _03779_ _03848_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09134__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ _03753_ _03758_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__xor2_4
XFILLER_0_98_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[16\] net878 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11229__B1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\] net770 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ net256 net2266 net474 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__mux2_1
XANTENNA__08645__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09842__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11521_ net913 _07117_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__nor2_1
XANTENNA__12247__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11452_ net334 net2566 net582 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
X_14240_ net1076 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10275__B _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ _04601_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__nor2_1
X_14171_ net1048 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ _06332_ _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15233__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] net991 _04276_ _04279_ vssd1
+ vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__or4b_4
XFILLER_0_46_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10334_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] net819 net766 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\]
+ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13053_ _02909_ _02947_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__xor2_1
X_10265_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\] net708 net696 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\]
+ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12004_ net238 net2352 net470 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XANTENNA__09373__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\] net816 net780 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16812_ net1366 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
XFILLER_0_79_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09125__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11834__B _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16743_ net1297 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
X_13955_ net1020 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ team_02_WB.instance_to_wrap.top.pc\[9\] _05635_ vssd1 vssd1 vccd1 vccd1 _02940_
+ sky130_fd_sc_hd__or2_1
X_16674_ net1229 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
X_13886_ net1021 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XANTENNA__10140__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__B2 team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15625_ clknet_leaf_29_wb_clk_i _02076_ _00583_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ _07369_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ clknet_leaf_55_wb_clk_i _02007_ _00514_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09833__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ _06266_ _05337_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14507_ net1013 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XANTENNA__12157__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ net267 net2726 net564 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__mux2_1
X_15487_ clknet_leaf_26_wb_clk_i _01938_ _00445_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12699_ _04592_ _06320_ _07325_ net826 vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 wbm_dat_i[12] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ net1139 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
Xinput21 wbm_dat_i[22] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 wbm_dat_i[3] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput43 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput54 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13393__B1 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput65 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
Xhold805 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ net1101 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
Xinput76 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold816 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16108_ clknet_leaf_64_wb_clk_i _02554_ _01066_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold827 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xinput98 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_1
Xhold838 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15726__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08930_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] net729 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16039_ clknet_leaf_15_wb_clk_i _02490_ _00997_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09364__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ net1564 _04558_ _04557_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07812_ _03670_ _03695_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__xnor2_1
X_08792_ net173 net953 net904 net1526 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09116__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15876__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _03599_ _03628_ _03631_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__nor3_1
XFILLER_0_135_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07674_ _03536_ _03563_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__xnor2_1
X_09413_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] net680 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12856__A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] net855 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a22o_1
XANTENNA__09824__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16699__1253 vssd1 vssd1 vccd1 vccd1 _16699__1253/HI net1253 sky130_fd_sc_hd__conb_1
XFILLER_0_48_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12067__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A _07215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08226_ _04089_ _04090_ _04082_ _04086_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a211o_1
XANTENNA__16501__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ _04008_ _04036_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10198__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08088_ _03946_ _03967_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10050_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\] net637 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12530__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14311__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09107__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ net1004 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
X_10952_ net399 _06590_ _06591_ _06592_ net416 vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__a221o_1
XANTENNA__10122__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13671_ net1152 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883_ _06100_ _06107_ net390 vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__mux2_1
XANTENNA__12766__A _05296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15410_ clknet_leaf_21_wb_clk_i _01861_ _00368_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _06473_ _07249_ _06482_ _06867_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__or4b_1
X_16390_ clknet_leaf_77_wb_clk_i _02821_ _01264_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15341_ clknet_leaf_23_wb_clk_i _01792_ _00299_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12553_ net308 net1768 net467 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10976__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11504_ _05839_ _05884_ _06007_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__nor3_1
X_15272_ clknet_leaf_56_wb_clk_i _01723_ _00230_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ net286 net2010 net481 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14223_ net1126 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11435_ net387 _07038_ net395 vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10189__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12705__S _07322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _06859_ _06976_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__nand2_1
X_14154_ net1036 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13105_ _02927_ _02933_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__xnor2_1
X_10317_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] net680 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\]
+ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__a221o_1
X_14085_ net1076 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
X_11297_ _06863_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15899__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ _02952_ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__xnor2_1
X_10248_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[2\] net785 _05902_ _05903_
+ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1130 net1133 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_4
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1141 net1142 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_4
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_4
XANTENNA__12440__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _05826_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nor2_8
Xfanout1163 net1165 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1174 net1185 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_4
Xfanout1185 net1205 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XANTENNA__15129__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1196 net1204 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_4
X_14987_ net1175 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16726_ net1280 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13938_ net1082 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08857__B2 net1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10664__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16657_ net1391 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_13869_ net1135 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15608_ clknet_leaf_123_wb_clk_i _02059_ _00566_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16588_ clknet_leaf_57_wb_clk_i net1407 _01461_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09806__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15539_ clknet_leaf_124_wb_clk_i _01990_ _00497_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14891__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _04722_ _04741_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ _03897_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10924__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold602 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold624 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold646 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold657 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[8\] net686 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08913_ _04584_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__or2_1
XANTENNA__09337__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09893_ _05550_ _05552_ _05554_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1302 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ net12 net950 _04555_ net2596 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a22o_1
XANTENNA__12350__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1313 team_02_WB.instance_to_wrap.top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 net2711
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1003_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1324 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1
+ net2722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1335 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 team_02_WB.instance_to_wrap.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net2744
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08775_ net1633 net956 net927 _04544_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XANTENNA__16054__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _03594_ _03615_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10104__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07657_ _03542_ _03543_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07588_ _03477_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09327_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] net722 _04501_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\]
+ _05002_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a221o_1
XANTENNA__09273__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09258_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\] net783 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08209_ _04089_ _04090_ _04073_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12525__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09189_ _04845_ _04866_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11220_ _05318_ _06183_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13109__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net909 _06295_ _06774_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10102_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\] net678 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__a22o_1
XANTENNA__09328__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ net396 _06466_ _06712_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10033_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[7\] net837 _05691_ _05693_
+ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a211o_1
X_14910_ net1170 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XANTENNA__12260__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ clknet_leaf_20_wb_clk_i _02341_ _00848_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A wbm_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ net1168 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14772_ net1181 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XANTENNA__08839__B2 team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11984_ net2156 net321 net534 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16511_ clknet_leaf_28_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[14\]
+ _01385_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13723_ net1058 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XANTENNA__09500__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10935_ net407 _06566_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11604__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16442_ clknet_leaf_90_wb_clk_i net1474 _01316_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ net1109 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
X_10866_ net413 net436 _06506_ _06510_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__a311o_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12605_ _06808_ _06870_ _07232_ _06842_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16373_ clknet_leaf_73_wb_clk_i net1691 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15571__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13585_ net1150 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10797_ net378 _06080_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15324_ clknet_leaf_63_wb_clk_i _01775_ _00282_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12536_ net252 net2263 net466 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15255_ clknet_leaf_118_wb_clk_i _01706_ _00213_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12467_ net239 net2203 net481 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XANTENNA__12435__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ net1070 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
X_11418_ net410 _06634_ _07023_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__o22a_1
XFILLER_0_50_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15186_ clknet_leaf_15_wb_clk_i _01637_ _00144_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12398_ net360 net2059 net492 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08775__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ net1063 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11349_ net393 _06762_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09319__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068_ net1039 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XANTENNA__16077__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16698__1252 vssd1 vssd1 vccd1 vccd1 _16698__1252/HI net1252 sky130_fd_sc_hd__conb_1
XANTENNA__12170__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _07385_ _07386_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10334__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ net72 net1593 net891 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07511_ net2084 net118 _00011_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ net1263 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08491_ _03420_ net961 vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nor2_1
XANTENNA__15914__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _04787_ _04789_ _04791_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or4_2
XFILLER_0_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12853__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09043_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\] net798 net790 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12345__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout309_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09558__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold410 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13965__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold454 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1120_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _04626_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
Xhold498 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout912 _04361_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_2
X_09945_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\] net811 _05606_ _05607_
+ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout923 _04555_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout580_A _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 _04355_ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_2
XANTENNA__12080__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout967 net970 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_2
X_09876_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\] net726 net708 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__a22o_1
XANTENNA__10325__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout978 team_02_WB.instance_to_wrap.top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ net978 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15444__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1110 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout989 team_02_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_8
Xhold1132 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ net31 net947 net921 net1702 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__o22a_1
XANTENNA__09730__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1143 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 net135 vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1176 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08758_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[13\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[13\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__mux2_2
Xhold1198 team_02_WB.instance_to_wrap.ramload\[14\] vssd1 vssd1 vccd1 vccd1 net2596
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _03597_ _03598_ _03558_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_71_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15594__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ net747 _04446_ _04455_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__and3_4
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10720_ _04763_ net373 vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ _06244_ _06302_ _06245_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] net930 net591 vssd1
+ vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13370_ _03216_ _03219_ _03239_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10800__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ net301 net1739 net502 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12255__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1154 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__inv_2
X_12252_ net270 net1714 net508 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08757__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A2 _06963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11203_ team_02_WB.instance_to_wrap.top.pc\[17\] _06336_ vssd1 vssd1 vccd1 vccd1
+ _06827_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12183_ net322 net1860 net519 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07873__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ net393 _06762_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15942_ clknet_leaf_12_wb_clk_i _02393_ _00900_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11065_ _06694_ _06697_ _06698_ team_02_WB.instance_to_wrap.top.aluOut\[22\] net459
+ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__o32a_4
XFILLER_0_120_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10316__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09182__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _05667_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10867__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15873_ clknet_leaf_3_wb_clk_i _02324_ _00831_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10867__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15937__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14824_ net1190 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ net1179 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11967_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ _04429_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10739__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10095__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ net1054 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10918_ _06046_ _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nor2_1
X_14686_ net1193 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11292__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11898_ net352 net2425 net544 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16425_ clknet_leaf_61_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[24\]
+ _01299_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13637_ net1087 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10849_ _06368_ _06375_ net363 vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ clknet_leaf_102_wb_clk_i _02789_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09788__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13568_ net1171 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08996__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ clknet_leaf_19_wb_clk_i _01758_ _00265_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15317__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12792__A1 _07410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12519_ net1775 net299 net476 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12165__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16287_ clknet_leaf_94_wb_clk_i _02720_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\] _03353_ _03337_ vssd1
+ vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ clknet_leaf_11_wb_clk_i _01689_ _00196_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ clknet_leaf_130_wb_clk_i _01620_ _00127_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09960__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ _03878_ _03846_ _03876_ _03879_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07971__B2 _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _04626_ team_02_WB.instance_to_wrap.top.DUT.read_data2\[14\] net592 vssd1
+ vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10307__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\] net708 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a22o_1
XANTENNA__09712__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08612_ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__inv_2
X_09592_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\] net864 net788 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11807__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ net80 net1563 net893 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10086__A2 _05725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08474_ net1525 net752 _04324_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1070_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout426_A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire609 _05112_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09779__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12075__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\] net665 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08739__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 team_02_WB.instance_to_wrap.top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1
+ net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold251 _02830_ vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_02_WB.START_ADDR_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07693__A team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10010__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09951__A2 _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 team_02_WB.instance_to_wrap.top.a1.row1\[1\] vssd1 vssd1 vccd1 vccd1 net1682
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_02_WB.START_ADDR_VAL_REG\[2\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout962_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout720 _04453_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
Xfanout731 _04448_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
X_09928_ _05581_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nor2_4
Xfanout742 _04324_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_4
Xfanout753 _04680_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_8
Xfanout764 _04675_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
Xfanout786 net788 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09703__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09859_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__inv_2
Xfanout797 net800 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12870_ _02903_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11821_ net300 net1991 net554 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07478__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ net1019 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
X_11752_ net269 net1838 net560 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10703_ _05134_ net368 vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14471_ net1153 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ net319 net1843 net571 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13015__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ clknet_leaf_36_wb_clk_i _02655_ _01167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input91_A wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _03304_ _03305_ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or3_1
X_10634_ _06264_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__or2_1
X_16697__1251 vssd1 vssd1 vccd1 vccd1 _16697__1251/HI net1251 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16141_ clknet_leaf_0_wb_clk_i net1500 _01099_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13353_ team_02_WB.instance_to_wrap.top.a1.row1\[2\] _03227_ _03238_ team_02_WB.instance_to_wrap.top.a1.row2\[34\]
+ _03256_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10565_ _04703_ _06215_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ net246 net1983 net500 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
X_16072_ clknet_leaf_85_wb_clk_i _02523_ _01030_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_13284_ _03181_ _03188_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10496_ _05442_ _06022_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15023_ net1189 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__inv_2
X_12235_ _04576_ _04578_ _07194_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__or3_4
XFILLER_0_62_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10001__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ net358 net1812 net522 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
XANTENNA__10741__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ team_02_WB.instance_to_wrap.top.pc\[20\] _06338_ vssd1 vssd1 vccd1 vccd1
+ _06747_ sky130_fd_sc_hd__nor2_1
X_12097_ net344 net2400 net524 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09155__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15925_ clknet_leaf_123_wb_clk_i _02376_ _00883_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11048_ net396 _06422_ _06681_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__o21a_1
Xinput8 wbm_dat_i[10] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15856_ clknet_leaf_34_wb_clk_i _02307_ _00814_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14807_ net1182 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15787_ clknet_leaf_21_wb_clk_i _02238_ _00745_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12999_ _02892_ _02893_ _02961_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10068__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ net1034 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14669_ net1043 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16408_ clknet_leaf_59_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[7\]
+ _01282_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08190_ _04039_ _04059_ _04056_ _04035_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__o211a_1
XANTENNA_wire596_A _05790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ clknet_leaf_99_wb_clk_i _02772_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08433__A2 _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10776__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10240__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09993__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09394__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09933__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__A team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07974_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] _03816_ _03827_ vssd1 vssd1
+ vccd1 vccd1 _03864_ sky130_fd_sc_hd__or3_1
XANTENNA__09146__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\] net806 net786 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\]
+ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12859__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09644_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[16\] net809 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[16\]
+ _05298_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08548__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09233__A _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\] net623 net619 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout543_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08526_ _04346_ _04347_ _04349_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or4_2
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10059__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08457_ net960 _04311_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout710_A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout808_A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15632__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08388_ _04248_ _04259_ _04251_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10350_ net398 _05882_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\] net786 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ net750 _05546_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__o21a_2
XANTENNA__15782__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09385__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ net267 net2126 net468 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
XANTENNA__09924__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _07200_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_8
Xfanout561 net563 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout572 _07191_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_8
Xfanout583 _04580_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
X_13971_ net1148 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12769__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _04577_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08966__B team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15710_ clknet_leaf_4_wb_clk_i _02161_ _00668_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12922_ _02900_ _02955_ _02901_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10298__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16690_ net1244 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08458__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ clknet_leaf_117_wb_clk_i _02092_ _00599_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09143__A _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ team_02_WB.instance_to_wrap.top.pc\[24\] _04629_ vssd1 vssd1 vccd1 vccd1
+ _02887_ sky130_fd_sc_hd__and2_1
XANTENNA__15162__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net246 net2196 net553 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ clknet_leaf_51_wb_clk_i _02023_ _00530_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08982__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12784_ _05836_ _05797_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14523_ net1048 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11735_ net594 _07188_ _07194_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08663__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11612__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454_ net1106 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11666_ net235 net2437 net574 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13405_ net1524 _04261_ net828 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
X_10617_ team_02_WB.instance_to_wrap.top.pc\[14\] _06268_ vssd1 vssd1 vccd1 vccd1
+ _06269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14385_ net1080 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
X_11597_ net236 net1862 net584 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
X_16124_ clknet_leaf_64_wb_clk_i _02570_ _01082_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10222__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ team_02_WB.instance_to_wrap.top.a1.row2\[24\] _03237_ _03238_ team_02_WB.instance_to_wrap.top.a1.row2\[32\]
+ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a221o_1
X_10548_ _06040_ _06199_ _06200_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16055_ clknet_leaf_118_wb_clk_i _02506_ _01013_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13267_ team_02_WB.instance_to_wrap.top.pad.keyCode\[7\] team_02_WB.instance_to_wrap.top.pad.keyCode\[6\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] team_02_WB.instance_to_wrap.top.pad.keyCode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__or4b_2
XANTENNA__12443__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10752__A _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ _04599_ _06130_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15006_ net1150 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
X_12218_ net325 net1867 net512 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__mux2_1
XANTENNA__09915__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ team_02_WB.START_ADDR_VAL_REG\[6\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net220 sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12149_ net315 net2220 net522 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09128__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15908_ clknet_leaf_53_wb_clk_i _02359_ _00866_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10289__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _03577_ _03578_ _03580_ _03571_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__o31a_2
X_15839_ clknet_leaf_26_wb_clk_i _02290_ _00797_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\] net701 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08892__A team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09300__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _04178_ _04184_ _04187_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09291_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] net729 net694 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08654__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08242_ _04100_ _04119_ _04102_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08173_ _04045_ _04049_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10213__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12353__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_112_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[1] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__09367__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__A2 _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 wbm_sel_o[1] sky130_fd_sc_hd__buf_2
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1200_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _03805_ _03824_ net262 _03796_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a31o_1
XANTENNA__15185__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16696__1250 vssd1 vssd1 vccd1 vccd1 _16696__1250/HI net1250 sky130_fd_sc_hd__conb_1
XANTENNA_fanout660_A _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__B net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12674__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _03748_ _03773_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_98_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09627_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[18\] net810 _05228_ _05229_
+ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ net988 team_02_WB.instance_to_wrap.wb.curr_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _04339_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08645__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12528__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\] net707 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ _05161_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XANTENNA__10988__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11520_ team_02_WB.instance_to_wrap.top.pc\[3\] team_02_WB.instance_to_wrap.top.pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11451_ team_02_WB.instance_to_wrap.top.aluOut\[7\] _07054_ _04582_ vssd1 vssd1 vccd1
+ vccd1 _07055_ sky130_fd_sc_hd__mux2_4
XFILLER_0_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ _04585_ _04597_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nand2_2
X_14170_ net1039 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11382_ team_02_WB.instance_to_wrap.top.pc\[9\] _06331_ team_02_WB.instance_to_wrap.top.pc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11668__A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ team_02_WB.instance_to_wrap.top.pc\[2\] net945 net942 _03125_ vssd1 vssd1
+ vccd1 vccd1 _01500_ sky130_fd_sc_hd__a22o_1
X_10333_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] net822 net862 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12263__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09358__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ team_02_WB.instance_to_wrap.top.pc\[14\] net944 net941 _03068_ vssd1 vssd1
+ vccd1 vccd1 _01512_ sky130_fd_sc_hd__a22o_1
X_10264_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] net712 net704 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a22o_1
XANTENNA__15528__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12003_ _04576_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__nand2_1
X_10195_ _05845_ _05847_ _05849_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16811_ net1365 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12499__A team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11607__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11468__A1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ net1093 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
X_16742_ net1296 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15678__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ _02917_ _02938_ _02915_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__o21a_1
X_16673_ net1228 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13885_ net1030 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12836_ _04804_ _06228_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__o21bai_1
X_15624_ clknet_leaf_110_wb_clk_i _02075_ _00582_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12968__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15555_ clknet_leaf_40_wb_clk_i _02006_ _00513_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12968__B2 _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12438__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12767_ _05337_ _06266_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__and2b_1
XANTENNA__10747__A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14506_ net1036 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11718_ net324 net2736 net564 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15486_ clknet_leaf_4_wb_clk_i _01937_ _00444_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12698_ _07324_ _07323_ _07322_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14437_ net1074 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
Xinput11 wbm_dat_i[13] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ net320 net2591 net575 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
Xinput22 wbm_dat_i[23] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput33 wbm_dat_i[4] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09597__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput44 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_14368_ net1076 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
Xinput66 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
Xinput77 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
Xhold806 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ clknet_leaf_64_wb_clk_i _02553_ _01065_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold817 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 team_02_WB.instance_to_wrap.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net2226
+ sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13319_ net985 team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] vssd1 vssd1 vccd1
+ vccd1 _03225_ sky130_fd_sc_hd__nand2b_1
Xhold839 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12173__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput99 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_1
XFILLER_0_64_1458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14299_ net1060 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XANTENNA__09349__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16038_ clknet_leaf_13_wb_clk_i _02489_ _00996_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08860_ net959 _04287_ _04299_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07811_ _03699_ _03700_ _03693_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ net1639 net953 net904 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[29\]
+ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07742_ _03599_ _03631_ _03632_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__or3b_1
XANTENNA__12202__A _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07673_ _03533_ _03536_ _03538_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09412_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\] net732 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07976__A2_N _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\] net824 net836 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[23\]
+ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a221o_1
XANTENNA__13081__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _04922_ _04931_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08277__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08225_ _04089_ _04090_ _04082_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _04015_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09052__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12083__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ _03946_ _03967_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_105_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11147__B1 team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15820__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net882 _04636_ _04648_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__and3_4
XFILLER_0_93_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09512__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ net383 _06443_ net393 vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15970__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13670_ net1141 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
X_10882_ net399 _06524_ _06525_ _06526_ net416 vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12621_ _06562_ _07248_ _06892_ _06545_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__or4b_1
XFILLER_0_13_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12258__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ clknet_leaf_53_wb_clk_i _01791_ _00298_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12552_ net301 net2198 net464 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09291__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11503_ net410 net449 _06739_ _07100_ _06630_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__o311a_1
XANTENNA__10830__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15271_ clknet_leaf_14_wb_clk_i _01722_ _00229_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12483_ net270 net2619 net480 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09579__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14222_ net1117 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_11434_ net383 _06960_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09043__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14153_ net1011 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
X_11365_ _05572_ _06174_ _06858_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13104_ team_02_WB.instance_to_wrap.top.pc\[5\] net945 net941 _03111_ vssd1 vssd1
+ vccd1 vccd1 _01503_ sky130_fd_sc_hd__a22o_1
X_10316_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] net664 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ net1142 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11296_ _06149_ _06178_ _06862_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__and3_1
X_13035_ _02904_ _02905_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\] net777 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\]
+ _05893_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__a221o_1
XANTENNA__14502__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1120 net1122 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_4
Xfanout1131 net1133 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_2
XFILLER_0_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09751__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1142 net1147 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
Xfanout1153 net1160 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_4
X_10178_ _05828_ _05830_ _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__or4_4
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_4
Xfanout1175 net1185 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_4
Xfanout1186 net1192 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
Xfanout1197 net1204 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_2
X_14986_ net1187 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
XANTENNA__09503__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16725_ net1279 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_89_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ net1028 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XANTENNA__08857__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10664__A2 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ net1004 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
X_16656_ net1390 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ clknet_leaf_117_wb_clk_i _02058_ _00565_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12819_ _05297_ _06263_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16587_ clknet_leaf_64_wb_clk_i net1440 _01460_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_13799_ net1152 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15538_ clknet_leaf_25_wb_clk_i _01989_ _00496_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09282__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15469_ clknet_leaf_23_wb_clk_i _01920_ _00427_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ _03866_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11800__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09034__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold603 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold614 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold658 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15843__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09961_ _05616_ _05618_ _05620_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__or4_2
XANTENNA__09990__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold669 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08912_ _04368_ net910 _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] net859 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[10\]
+ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__a221o_1
XANTENNA__10940__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net13 net948 net922 net1647 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1303 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08410__A _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1314 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 team_02_WB.instance_to_wrap.top.a1.row1\[16\] vssd1 vssd1 vccd1 vccd1 net2723
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1336 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1347 team_02_WB.instance_to_wrap.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net2745
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08774_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[5\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[5\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__mux2_2
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _03581_ _03604_ _03594_ _03590_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__A team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1198_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07656_ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] _03476_ _03510_ _03545_ _03546_
+ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o32a_2
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15223__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08556__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12078__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_A _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _03446_ _03474_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09326_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\] net678 net663 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\]
+ _04996_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09273__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15373__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[25\] net823 net776 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08208_ team_02_WB.instance_to_wrap.top.a1.row2\[32\] net936 net919 _04091_ vssd1
+ vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09025__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08139_ _03988_ _04011_ _04014_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nand4_1
XFILLER_0_47_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11150_ _06255_ net743 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] net443
+ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a221o_1
XANTENNA__09981__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10101_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\] net734 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\]
+ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11081_ _06713_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__inv_2
XANTENNA__12541__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\] net785 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[7\]
+ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a221o_1
XANTENNA__08000__A3 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ net1168 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A wbm_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1199 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
X_11983_ net2401 net316 net533 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08839__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12777__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ net1058 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
X_16510_ clknet_leaf_6_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[13\]
+ _01384_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10934_ net408 _06576_ _06573_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ net1118 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
X_16441_ clknet_leaf_89_wb_clk_i net1480 _01315_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10865_ _04824_ net430 _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__a21o_1
XANTENNA__15716__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ _06894_ _06927_ _06939_ _07231_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__nand4_1
X_16372_ clknet_leaf_73_wb_clk_i _02803_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ net1150 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09264__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10796_ _06443_ _06444_ net387 vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15323_ clknet_leaf_119_wb_clk_i _01774_ _00281_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12535_ net249 net2652 net466 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15254_ clknet_leaf_109_wb_clk_i _01705_ _00212_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12466_ _07199_ _07214_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15866__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14205_ net1080 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_11417_ net398 _06849_ net410 vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15185_ clknet_leaf_19_wb_clk_i _01636_ _00143_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12397_ net352 net2110 net492 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10031__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B2 _04544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14136_ net1107 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11348_ _06872_ _06960_ net383 vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10582__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net1144 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XANTENNA__12451__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _06680_ _06897_ net394 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10760__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13018_ net232 _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15246__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14969_ net1002 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07510_ team_02_WB.instance_to_wrap.top.pad.count\[0\] team_02_WB.instance_to_wrap.top.pad.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16708_ net1262 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
X_08490_ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] _04275_ _04326_ vssd1 vssd1
+ vccd1 vccd1 _04327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15396__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16639_ net1210 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09996__A _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\] net684 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[28\]
+ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09042_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[30\] net809 net805 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\]
+ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a221o_1
XANTENNA__10270__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold400 team_02_WB.instance_to_wrap.top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 net1798
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold411 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold422 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09963__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold444 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10573__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16021__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold488 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\] net880 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ _05596_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a221o_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12361__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold499 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1113_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 net927 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net938 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09715__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout946 _07363_ vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_2
XANTENNA_input9_A wbm_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_2
X_09875_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\] net682 net661 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\]
+ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a221o_1
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
Xhold1100 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A _07191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 team_02_WB.instance_to_wrap.top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1
+ net979 sky130_fd_sc_hd__clkbuf_4
Xhold1111 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ team_02_WB.instance_to_wrap.busy_o net949 team_02_WB.instance_to_wrap.wb.prev_BUSY_O
+ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1133 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 team_02_WB.START_ADDR_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\] vssd1 vssd1 vccd1 vccd1
+ net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net1617 net957 net926 _04535_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1177 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11705__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] net654 net650 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ _04482_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a221o_1
XANTENNA__09494__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07639_ _03492_ _03525_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10650_ team_02_WB.instance_to_wrap.top.pc\[22\] _06246_ _06301_ vssd1 vssd1 vccd1
+ vccd1 _06302_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15889__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09246__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11589__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09309_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[24\] net782 net758 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[24\]
+ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ team_02_WB.instance_to_wrap.top.pc\[27\] _06231_ vssd1 vssd1 vccd1 vccd1
+ _06233_ sky130_fd_sc_hd__or2_1
XANTENNA__12536__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14317__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10261__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ net292 net2633 net501 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ net323 net2669 net508 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10013__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ net442 _06808_ _06810_ _06826_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[17\]
+ sky130_fd_sc_hd__a211o_2
XANTENNA__08757__B2 _04535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net315 net2148 net517 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11133_ _06649_ _06761_ net382 vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12271__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09706__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16514__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11064_ _06246_ net743 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] net443
+ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__a221o_1
X_15941_ clknet_leaf_128_wb_clk_i _02392_ _00899_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _05669_ _05671_ _05673_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ clknet_leaf_9_wb_clk_i _02323_ _00830_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14823_ net1188 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11615__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ net233 net1744 net538 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
X_14754_ net1178 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09485__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__A1 team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ net1024 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
X_10917_ _04913_ _06045_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__nor2_1
X_14685_ net1194 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08693__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ net354 net2606 net547 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16424_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[23\]
+ _01298_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_13636_ net1093 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848_ _06490_ _06494_ net404 vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16355_ clknet_leaf_102_wb_clk_i _02788_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13567_ net1172 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__inv_2
XANTENNA__12446__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ net439 _06410_ _06427_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15306_ clknet_leaf_44_wb_clk_i _01757_ _00264_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12518_ net1814 net294 net476 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16286_ clknet_leaf_95_wb_clk_i _02719_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13498_ _03353_ net873 _03352_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16044__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ clknet_leaf_125_wb_clk_i _01688_ _00195_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12449_ net324 net2504 net484 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10004__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15168_ clknet_leaf_8_wb_clk_i _01619_ _00126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14119_ net1153 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12181__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ _03878_ _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nand2b_1
X_15099_ clknet_leaf_119_wb_clk_i _01550_ _00057_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\] net685 net664 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ _03396_ _04406_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__or3_2
XFILLER_0_136_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\] net819 net836 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08542_ net81 net1636 net892 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__A1 team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08473_ team_02_WB.instance_to_wrap.top.a1.state\[2\] net752 vssd1 vssd1 vccd1 vccd1
+ _04324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12356__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10243__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\] net736 _04708_ vssd1
+ vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07974__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15411__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold230 team_02_WB.instance_to_wrap.top.a1.row1\[112\] vssd1 vssd1 vccd1 vccd1 net1628
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 net174 vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A _04468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold263 team_02_WB.START_ADDR_VAL_REG\[4\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12091__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 team_02_WB.instance_to_wrap.top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1 net1672
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 team_02_WB.instance_to_wrap.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net1683
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold296 team_02_WB.START_ADDR_VAL_REG\[25\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _04458_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_8
Xfanout721 _04453_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
Xfanout732 _04447_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09927_ _05583_ _05585_ _05587_ _05589_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__or4_2
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout955_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 _04680_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
Xfanout765 _04674_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 _04671_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
X_09858_ _05503_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__nand2_1
Xfanout798 net800 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_4
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08809_ net155 net954 net905 net1545 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
X_09789_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[12\] net661 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\]
+ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11820_ net291 net2482 net552 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09467__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11751_ net324 net2404 net560 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XANTENNA__08675__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ _05175_ net372 vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14470_ net1092 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
X_11682_ net317 net2602 net570 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13421_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[17\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16067__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10633_ team_02_WB.instance_to_wrap.top.pc\[16\] _06263_ vssd1 vssd1 vccd1 vccd1
+ _06285_ sky130_fd_sc_hd__nor2_1
XANTENNA__13038__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12266__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10234__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16140_ clknet_leaf_129_wb_clk_i net1502 _01098_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dfrtp_1
X_13352_ net896 _03244_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__nand2_1
XANTENNA_input84_A wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _04703_ _06215_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ net242 net2559 net500 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XANTENNA__13886__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16071_ clknet_leaf_14_wb_clk_i _02522_ _01029_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13283_ net1638 _03174_ _03187_ _03194_ net995 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__inv_2
XANTENNA__12790__A _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15022_ net1190 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ net233 net2179 net514 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16627__1206 vssd1 vssd1 vccd1 vccd1 _16627__1206/HI net1206 sky130_fd_sc_hd__conb_1
X_12165_ net353 net2028 net520 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net440 _06729_ _06730_ net427 _06746_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[20\]
+ sky130_fd_sc_hd__o221ai_4
XFILLER_0_21_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12096_ net348 net2335 net526 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
X_15924_ clknet_leaf_46_wb_clk_i _02375_ _00882_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11047_ net401 _06417_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a21bo_1
Xinput9 wbm_dat_i[11] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_1
X_15855_ clknet_leaf_31_wb_clk_i _02306_ _00813_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14806_ net1201 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15786_ clknet_leaf_46_wb_clk_i _02237_ _00744_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09458__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12998_ team_02_WB.instance_to_wrap.top.pc\[23\] net943 net942 _03023_ vssd1 vssd1
+ vccd1 vccd1 _01521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14737_ net1008 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
X_11949_ net320 net2145 net539 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ net1033 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16407_ clknet_leaf_75_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[6\]
+ _01281_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12176__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ net1127 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14599_ net1178 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15434__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10916__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16338_ clknet_leaf_99_wb_clk_i _02771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09091__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16269_ clknet_leaf_79_wb_clk_i _02702_ _01221_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ _03861_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nand2_1
X_09712_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] net782 net767 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09697__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] net865 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\]
+ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout271_A _06674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout369_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09574_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\] net635 net631 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a22o_1
XANTENNA__09449__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ _04350_ _04351_ _04352_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__or4_1
XANTENNA__11256__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout536_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08456_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[3\] net917 vssd1 vssd1 vccd1
+ vccd1 _04312_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _04249_ _04250_ _04252_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12086__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09621__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15927__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09008_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net857 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10280_ _04505_ _04507_ _05886_ net462 net740 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout540 _07202_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_6
Xfanout551 _07200_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11599__C_N team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_8
Xfanout573 _07191_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_4
X_13970_ net1084 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XANTENNA__12141__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout584 _04580_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_6
X_12921_ team_02_WB.instance_to_wrap.top.pc\[17\] _06263_ _02954_ vssd1 vssd1 vccd1
+ vccd1 _02955_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15307__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15640_ clknet_leaf_122_wb_clk_i _02091_ _00598_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12852_ team_02_WB.instance_to_wrap.top.pc\[25\] _06241_ vssd1 vssd1 vccd1 vccd1
+ _02886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net242 net2268 net553 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ clknet_leaf_125_wb_clk_i _02022_ _00529_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12783_ _05768_ _05771_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__and2b_1
XANTENNA__12785__A _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08982__B _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14522_ net1046 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11734_ net235 net2262 net567 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ net1121 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
X_11665_ net359 net2016 net574 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ net750 _05841_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__o21a_2
X_13404_ net1505 _04263_ net828 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
XANTENNA__09073__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14384_ net1017 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
XANTENNA_output190_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11596_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[0\] _07185_ vssd1 vssd1 vccd1
+ vccd1 _07186_ sky130_fd_sc_hd__a21o_2
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09612__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ clknet_leaf_62_wb_clk_i _02569_ _01081_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13335_ team_02_WB.instance_to_wrap.top.a1.row1\[120\] _03239_ _03240_ team_02_WB.instance_to_wrap.top.a1.row2\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ _05012_ _05031_ _06145_ _06196_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08820__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13157__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ team_02_WB.instance_to_wrap.top.pad.keyCode\[2\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__or4b_2
X_16054_ clknet_leaf_111_wb_clk_i _02505_ _01012_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ _04599_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and2_1
X_12217_ net321 net2091 net515 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__mux2_1
X_15005_ net1147 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13197_ team_02_WB.START_ADDR_VAL_REG\[5\] net997 net933 vssd1 vssd1 vccd1 vccd1
+ net219 sky130_fd_sc_hd__a21o_1
X_16789__1343 vssd1 vssd1 vccd1 vccd1 _16789__1343/HI net1343 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12148_ net304 net2616 net523 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net279 net1875 net524 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XANTENNA__09679__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ clknet_leaf_41_wb_clk_i _02358_ _00865_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12780__A_N _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15838_ clknet_leaf_4_wb_clk_i _02289_ _00796_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15769_ clknet_leaf_107_wb_clk_i _02220_ _00727_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08892__B _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11803__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08310_ _04184_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16745__1299 vssd1 vssd1 vccd1 vccd1 _16745__1299/HI net1299 sky130_fd_sc_hd__conb_1
X_09290_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] net684 net662 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\]
+ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08241_ _04121_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08172_ _04019_ _04044_ _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__or4_4
XANTENNA__09064__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09603__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08811__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_99_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__clkbuf_4
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_112_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[30] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 wbm_sel_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__12910__A2 _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_10_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout486_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03842_ _03845_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07887_ _03707_ _03777_ _03774_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout653_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ _05286_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nor2_8
X_09557_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] net813 net798 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout918_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ net1766 _04338_ _04325_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
X_09488_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\] net631 net623 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a22o_1
XANTENNA__09842__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08439_ team_02_WB.instance_to_wrap.top.a1.data\[7\] net915 vssd1 vssd1 vccd1 vccd1
+ _04299_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11450_ team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] net887 net907 team_02_WB.instance_to_wrap.top.pc\[7\]
+ _07053_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09055__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10401_ _04703_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08802__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12544__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _05571_ _06135_ _06991_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[10\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120_ team_02_WB.instance_to_wrap.top.pc\[2\] net227 _03124_ vssd1 vssd1 vccd1
+ vccd1 _03125_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] net860 net756 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13051_ net889 _07439_ _03064_ _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__o31ai_1
X_10263_ _05911_ _05913_ _05915_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__or4_1
X_12002_ _07188_ _07205_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__nor2_1
XANTENNA__12901__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] net812 net764 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\]
+ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16810_ net1364 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_2
Xfanout381 _05955_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_2
Xfanout392 _05908_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_2
X_16741_ net1295 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XFILLER_0_96_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13953_ net1102 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12904_ _02920_ _02937_ _02918_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__o21a_1
X_16672_ net1227 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
X_13884_ net1102 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XANTENNA__10140__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15623_ clknet_leaf_14_wb_clk_i _02074_ _00581_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12835_ _07371_ _02868_ _07370_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11623__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15554_ clknet_leaf_47_wb_clk_i _02005_ _00512_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12766_ _05296_ _06263_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09833__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10747__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14505_ net1028 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11717_ net320 net1956 net567 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12697_ _04435_ _04591_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__or2_1
X_15485_ clknet_leaf_113_wb_clk_i _01936_ _00443_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ net317 net2676 net574 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XANTENNA__09046__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14436_ net1094 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
Xinput12 wbm_dat_i[14] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 wbm_dat_i[24] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 wbm_dat_i[5] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput45 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14367_ net1132 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XANTENNA__12454__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ net359 net2191 net583 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
Xinput56 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xhold807 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16106_ clknet_leaf_63_wb_clk_i _02552_ _01064_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput78 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10600__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput89 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
Xhold818 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ team_02_WB.instance_to_wrap.top.a1.row1\[16\] _03222_ _03223_ team_02_WB.instance_to_wrap.top.a1.row1\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a22o_1
Xhold829 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ net1039 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
X_16037_ clknet_leaf_125_wb_clk_i _02488_ _00995_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13249_ net2747 net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[22\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_21_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07810_ _03699_ _03700_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nand2_2
X_08790_ net1656 net953 net904 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XANTENNA__15622__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _03595_ _03615_ _03616_ _03593_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09521__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ _03533_ _03538_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] net712 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15772__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09342_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\] net808 net784 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__a22o_1
XANTENNA__09285__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09824__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09273_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[25\] net593 vssd1
+ vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08224_ _04069_ _04101_ _04104_ _04080_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08155_ _04011_ _04014_ _04024_ _04032_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__and4_2
XANTENNA__12364__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10198__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08086_ _03903_ _03945_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__or2_1
XANTENNA__08143__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15152__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11147__A1 team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout770_A _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16510__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08988_ net883 _04641_ _04648_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__and3_4
X_07939_ _03828_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10950_ net382 _06442_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__nand2_1
XANTENNA__10122__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] net716 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[16\]
+ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10881_ net387 _06084_ net394 vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__o21a_1
XANTENNA__12539__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input101_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ _06589_ _06666_ _07247_ _06914_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__or4b_1
XFILLER_0_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16788__1342 vssd1 vssd1 vccd1 vccd1 _16788__1342/HI net1342 sky130_fd_sc_hd__conb_1
XFILLER_0_136_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12551_ net291 net2342 net464 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ net410 _06739_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__nor2_1
XANTENNA__10830__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08752__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12482_ net325 net1794 net480 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__mux2_1
X_15270_ clknet_leaf_12_wb_clk_i _01721_ _00228_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12782__B _05725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14221_ net1132 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
X_11433_ _07001_ _07037_ net377 vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__mux2_1
XANTENNA__12274__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10189__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11386__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__B2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14152_ net1099 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
X_11364_ net310 net2358 net585 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13894__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ _07422_ _03108_ _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__o21ai_1
X_10315_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\] net674 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\]
+ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a221o_1
X_14083_ net1070 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ net283 net2462 net583 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13034_ _07366_ _03053_ team_02_WB.instance_to_wrap.top.pc\[17\] net943 vssd1 vssd1
+ vccd1 vccd1 _01515_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15645__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10246_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] net817 net814 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09200__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16744__1298 vssd1 vssd1 vccd1 vccd1 _16744__1298/HI net1298 sky130_fd_sc_hd__conb_1
Xfanout1110 net1113 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11618__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_4
X_10177_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\] net704 net701 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__a221o_1
Xfanout1143 net1145 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 net1160 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1169 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1176 net1184 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
Xfanout1187 net1192 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
X_14985_ net1191 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__inv_2
Xfanout1198 net1202 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_4
XANTENNA__15795__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16724_ net1278 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13936_ net1018 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16655_ net1389 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__12449__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ net1026 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
X_15606_ clknet_leaf_110_wb_clk_i _02057_ _00564_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12818_ _07390_ _07441_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__and2_1
X_16586_ clknet_leaf_65_wb_clk_i net1461 _01459_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09267__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13798_ net1139 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XANTENNA__09806__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15537_ clknet_leaf_18_wb_clk_i _01988_ _00495_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12749_ _04888_ _06234_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15468_ clknet_leaf_22_wb_clk_i _01919_ _00426_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15175__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ net1103 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16420__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12184__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15399_ clknet_leaf_14_wb_clk_i _01850_ _00357_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold604 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09059__A _04722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold615 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold626 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold637 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold648 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09960_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net714 net690 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__a221o_1
Xhold659 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12326__A0 _07055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08898__A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08911_ _04368_ _04593_ _04594_ _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__or4b_2
XANTENNA__16570__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[10\] net811 net842 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08842_ net14 net948 net922 net1836 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__o22a_1
Xhold1304 net129 vssd1 vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 team_02_WB.instance_to_wrap.top.a1.row1\[60\] vssd1 vssd1 vccd1 vccd1 net2713
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] vssd1
+ vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ net1729 net956 net925 _04543_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
Xhold1348 team_02_WB.instance_to_wrap.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net2746
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07724_ _03581_ _03604_ _03590_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10104__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__A _05175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _03511_ _03512_ _03537_ _03509_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__o211a_1
XANTENNA__12359__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_A _07153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09258__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07586_ team_02_WB.instance_to_wrap.top.a1.dataIn\[18\] _03474_ _03475_ vssd1 vssd1
+ vccd1 vccd1 _03477_ sky130_fd_sc_hd__or3_1
X_09325_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[23\] net711 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11065__B1 team_02_WB.instance_to_wrap.top.aluOut\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15518__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09256_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\] net868 net795 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12094__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09187_ _04845_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15668__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _03982_ _04017_ _04019_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__or3_2
XFILLER_0_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09430__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10040__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ _03925_ _03952_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[5\] net690 net670 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11080_ net396 _06462_ _06712_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__o21a_1
X_10031_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[7\] net861 net841 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ net1199 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
X_11982_ net1900 net303 net534 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XANTENNA__12777__B _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ net1058 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
X_10933_ _06574_ _06575_ net405 vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__mux2_1
XANTENNA__12269__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16440_ clknet_leaf_99_wb_clk_i net1468 _01314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13652_ net1038 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ _04826_ net452 net445 _04825_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__a22o_1
XANTENNA__13045__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _06958_ _06999_ _07230_ _06978_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16371_ clknet_leaf_74_wb_clk_i net1463 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.debounce_dly
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12991__A_N _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13583_ net1150 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
X_10795_ _06063_ _06089_ net363 vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15322_ clknet_leaf_120_wb_clk_i _01773_ _00280_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12534_ net245 net2309 net466 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15253_ clknet_leaf_124_wb_clk_i _01704_ _00211_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12465_ net233 net2129 net486 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12556__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14204_ net1085 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_11416_ net404 _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__nor2_1
X_15184_ clknet_leaf_39_wb_clk_i _01635_ _00142_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12396_ net355 net1986 net495 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09421__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14135_ net1112 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
X_11347_ _06916_ _06959_ net376 vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11278_ _06790_ _06896_ net385 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14066_ net1084 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10229_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] _04367_ _04426_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a22o_1
X_13017_ _02899_ _02956_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10334__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[8\] vssd1 vssd1 vccd1 vccd1
+ net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09488__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14968_ net1008 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16707_ net1261 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_72_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13919_ net1130 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12179__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14899_ net1171 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16638_ net1209 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16569_ clknet_leaf_99_wb_clk_i net1420 _01442_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09110_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] net697 net633 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11811__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09660__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] net866 net773 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09412__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold401 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold434 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15960__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09943_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[9\] net822 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
Xhold489 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout903 net905 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout914 _04361_ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_2
XFILLER_0_0_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16787__1341 vssd1 vssd1 vccd1 vccd1 _16787__1341/HI net1341 sky130_fd_sc_hd__conb_1
XANTENNA_fanout399_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
X_09874_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[10\] net730 net670 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a22o_1
Xfanout958 _04340_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
XANTENNA__10325__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_2
Xhold1101 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09191__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ team_02_WB.instance_to_wrap.busy_o team_02_WB.instance_to_wrap.wb.prev_BUSY_O
+ net948 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__and3b_2
Xhold1123 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1134 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _07195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 team_02_WB.instance_to_wrap.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net2554
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[14\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[14\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_1
Xhold1178 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
X_07707_ _03555_ _03572_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12089__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout733_A _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ net748 _04445_ _04449_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__and3_1
XANTENNA__15340__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07638_ _03494_ _03527_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07569_ _03458_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16743__1297 vssd1 vssd1 vccd1 vccd1 _16743__1297/HI net1297 sky130_fd_sc_hd__conb_1
XANTENNA__11721__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\] net850 net830 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10580_ team_02_WB.instance_to_wrap.top.pc\[27\] _06231_ vssd1 vssd1 vccd1 vccd1
+ _06232_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09651__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09239_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[25\] net700 net677 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a22o_1
XANTENNA__13221__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12538__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ net320 net1915 net511 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09403__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ net438 _06814_ _06823_ net449 _06825_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__a221o_1
XANTENNA__08757__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12181_ net305 net1793 net519 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12552__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _06708_ _06760_ net376 vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold990 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15940_ clknet_leaf_54_wb_clk_i _02391_ _00898_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ net912 _06696_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10316__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[7\] net708 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ _05674_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09182__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ clknet_leaf_27_wb_clk_i _02322_ _00829_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12788__A _07410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822_ net1188 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14753_ net1181 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11965_ net360 net2057 net536 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ net1100 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ _06307_ _06558_ net909 vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14684_ net1196 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09890__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net343 net2534 net545 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16423_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[22\]
+ _01297_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ net1068 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _06491_ _06493_ net391 vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11631__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16354_ clknet_leaf_102_wb_clk_i _02787_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13566_ net1172 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10788__C1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09642__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _04742_ net431 net447 _04743_ _06428_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15305_ clknet_leaf_29_wb_clk_i _01756_ _00263_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08996__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12517_ net2613 net284 net478 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
X_16285_ clknet_leaf_101_wb_clk_i _02718_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15983__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ _03134_ _03348_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15236_ clknet_leaf_19_wb_clk_i _01687_ _00194_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ net322 net1811 net487 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12462__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ clknet_leaf_27_wb_clk_i _01618_ _00125_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12379_ net298 net1929 net492 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15213__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16339__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ net1140 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15098_ clknet_leaf_121_wb_clk_i _01549_ _00056_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14049_ net1100 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10307__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15363__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11806__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ net975 net974 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__nand2b_1
X_09590_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net808 net772 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\]
+ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08541_ net82 net1606 net893 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11107__A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ _03420_ _04284_ net1675 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a21o_1
XANTENNA__13009__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13009__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11541__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09633__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13041__B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout314_A _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\] net680 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12880__B _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_02_WB.instance_to_wrap.top.pc\[2\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12372__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 net123 vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _02608_ vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold253 team_02_WB.instance_to_wrap.top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1 net1651
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 net136 vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold275 team_02_WB.instance_to_wrap.ramload\[1\] vssd1 vssd1 vccd1 vccd1 net1673
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
XFILLER_0_1_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold286 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 team_02_WB.START_ADDR_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15706__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13992__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout711 _04458_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
X_09926_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[9\] net657 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[9\]
+ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a221o_1
Xfanout722 _04453_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_6
Xfanout733 _04447_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 _06323_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
Xfanout755 _04680_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_8
Xfanout766 _04674_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_A _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[11\] net592 vssd1
+ vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__o21ai_4
Xfanout777 _04670_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
Xfanout788 _04665_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08372__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08808_ net156 net952 net902 net1519 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] net734 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a22o_1
XANTENNA__15856__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16674__1229 vssd1 vssd1 vccd1 vccd1 _16674__1229/HI net1229 sky130_fd_sc_hd__conb_1
X_08739_ net2552 net955 net924 _04526_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
XANTENNA__13216__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ net320 net2308 net563 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09872__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _06350_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12547__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ net305 net2436 net571 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__mux2_1
XANTENNA__11451__S _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__A team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__or4bb_1
X_10632_ team_02_WB.instance_to_wrap.top.pc\[15\] _06266_ _06283_ vssd1 vssd1 vccd1
+ vccd1 _06284_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09624__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13351_ team_02_WB.instance_to_wrap.top.a1.row1\[10\] _03223_ _03237_ team_02_WB.instance_to_wrap.top.a1.row2\[26\]
+ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a22o_1
X_10563_ _04702_ _06215_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08045__B _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15236__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ net237 net2740 net500 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070_ clknet_leaf_14_wb_clk_i _02521_ _01028_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input77_A wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13282_ _03189_ _03192_ _03193_ _03190_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or4b_1
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _05523_ _05524_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__nor2_2
XANTENNA__08760__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12790__B _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ net1189 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__inv_2
XANTENNA__12282__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ net359 net2483 net512 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__mux2_1
XANTENNA__10591__A team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12164_ net355 net2021 net523 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15386__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net439 _06734_ _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ net339 net2412 net526 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09155__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15923_ clknet_leaf_125_wb_clk_i _02374_ _00881_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11046_ net397 _06680_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__nand2_1
XANTENNA__11626__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15854_ clknet_leaf_33_wb_clk_i _02305_ _00812_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10170__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14805_ net1199 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15785_ clknet_leaf_32_wb_clk_i _02236_ _00743_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12997_ net229 _03019_ _03022_ _04362_ _03020_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12998__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14736_ net1033 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
X_11948_ net317 net2227 net537 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
XANTENNA__09863__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14667_ net1042 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12457__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14238__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ net289 net1877 net544 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16406_ clknet_leaf_76_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[5\]
+ _01280_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ net1078 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16786__1340 vssd1 vssd1 vccd1 vccd1 _16786__1340/HI net1340 sky130_fd_sc_hd__conb_1
XANTENNA__09615__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14598_ net1178 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11485__A2_N net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16337_ clknet_leaf_100_wb_clk_i _02770_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13549_ net1668 _03385_ net884 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11973__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16161__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16268_ clknet_leaf_92_wb_clk_i _02701_ _01220_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ clknet_leaf_3_wb_clk_i _01670_ _00177_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15729__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_81_wb_clk_i _02644_ _01156_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09394__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07972_ _03835_ _03860_ _03839_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09146__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16742__1296 vssd1 vssd1 vccd1 vccd1 _16742__1296/HI net1296 sky130_fd_sc_hd__conb_1
X_09711_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\] net849 net785 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a22o_1
XANTENNA__10161__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[17\] net666 _05243_ vssd1
+ vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__a21o_1
X_08524_ net56 net55 net58 net57 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09854__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07969__B _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ team_02_WB.instance_to_wrap.top.a1.data\[3\] net915 vssd1 vssd1 vccd1 vccd1
+ _04311_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout431_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1173_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08409__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08386_ _04250_ _04254_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13987__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _04685_ _04687_ _04689_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16513__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07526__A_N team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09385__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 _07202_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09909_ _05570_ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nor2_2
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_6
Xfanout563 _07196_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_8
Xfanout574 _07191_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_6
Xfanout585 _04580_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
X_12920_ _02902_ _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__and2b_1
XANTENNA__13227__A net1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12851_ team_02_WB.instance_to_wrap.top.pc\[26\] _06238_ vssd1 vssd1 vccd1 vccd1
+ _02885_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ net237 net2409 net552 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ clknet_leaf_25_wb_clk_i _02021_ _00528_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09845__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12782_ _05722_ _05725_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12785__B _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14521_ net1064 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09440__A _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net358 net2105 net564 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12277__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ net1034 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11664_ net352 net2367 net572 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13403_ net1489 _04265_ net828 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
X_10615_ net929 _05886_ _06220_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ net1123 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11595_ team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] net887 _07168_ team_02_WB.instance_to_wrap.top.pc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__a22o_1
X_16122_ clknet_leaf_63_wb_clk_i _02568_ _01080_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ _03209_ _03233_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10546_ _05053_ _05072_ _05075_ _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ clknet_leaf_114_wb_clk_i _02504_ _01011_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13265_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] _03177_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.lcd_en sky130_fd_sc_hd__a21oi_1
X_10477_ _04585_ _04596_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__nor2_1
X_15004_ net1188 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12216_ net315 net2476 net513 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ team_02_WB.START_ADDR_VAL_REG\[4\] _04356_ vssd1 vssd1 vccd1 vccd1 net218
+ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12147_ net295 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] net520 vssd1
+ vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09128__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12078_ net273 net2051 net526 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_15906_ clknet_leaf_47_wb_clk_i _02357_ _00864_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11029_ _06040_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__xor2_1
XANTENNA__10143__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15837_ clknet_leaf_114_wb_clk_i _02288_ _00795_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15768_ clknet_leaf_122_wb_clk_i _02219_ _00726_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09836__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16527__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__A1_N _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11643__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14719_ net1035 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12187__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15699_ clknet_leaf_124_wb_clk_i _02150_ _00657_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_08240_ _04101_ _04119_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__xnor2_2
XANTENNA_hold85_A team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08171_ _04044_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16673__1228 vssd1 vssd1 vccd1 vccd1 _16673__1228/HI net1228 sky130_fd_sc_hd__conb_1
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[11] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13022__A1_N _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09367__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[31] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 wbm_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__09119__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ _03809_ _03843_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout479_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ _03737_ _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _05288_ _05290_ _05292_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__or4_2
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout646_A _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] net863 net858 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a22o_1
XANTENNA__09827__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ _02861_ _04326_ _04334_ team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ _04279_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__o221a_1
XANTENNA__12097__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16508__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\] net695 net663 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ net1826 net827 _03423_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08369_ _04234_ _04235_ _04238_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a211o_1
X_10400_ _04744_ _06052_ _04742_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ net426 _06977_ _06978_ _04605_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[0\] net856 net836 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10262_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] net676 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a221o_1
XANTENNA__09358__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13050_ net230 _03066_ net227 _06908_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__o2bb2a_1
X_12001_ net2043 net235 net534 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
X_10193_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[3\] net864 net776 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a22o_1
XANTENNA__12560__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
Xfanout371 _05998_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_2
X_16740_ net1294 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
X_13952_ net1075 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10125__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12903_ _02923_ _02936_ _02921_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o21a_1
X_16671_ net1226 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__09530__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ net1047 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
XANTENNA__11904__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15622_ clknet_leaf_3_wb_clk_i _02073_ _00580_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12834_ _07372_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__A0 _07055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15553_ clknet_leaf_1_wb_clk_i _02004_ _00511_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16418__D team_02_WB.instance_to_wrap.top.ru.dmmload_co\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ _05257_ _06260_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11205__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14504_ net1083 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
X_11716_ net317 net2710 net566 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15484_ clknet_leaf_50_wb_clk_i _01935_ _00442_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12696_ _04435_ _06325_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14435_ net1068 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16741__1295 vssd1 vssd1 vccd1 vccd1 _16741__1295/HI net1295 sky130_fd_sc_hd__conb_1
X_11647_ net305 net2662 net575 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 wbm_dat_i[15] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 wbm_dat_i[25] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09597__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 wbm_dat_i[6] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
X_14366_ net1021 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
Xinput46 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_11578_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[1\] _07169_ vssd1 vssd1 vccd1
+ vccd1 _07170_ sky130_fd_sc_hd__a21o_2
XFILLER_0_29_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput57 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput68 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_1
X_16105_ clknet_leaf_70_wb_clk_i _02551_ _01063_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold808 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13317_ net986 net987 _03221_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold819 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ _06152_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput79 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
X_14297_ net1061 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ clknet_leaf_19_wb_clk_i _02487_ _00994_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09349__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ net1689 net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12470__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13179_ _02783_ _03161_ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07740_ _03597_ _03625_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10116__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _03529_ _03561_ _03556_ _03532_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15917__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] net728 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11616__A0 _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[23\] net859 net787 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ _05017_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09272_ _04941_ _04950_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[25\]
+ sky130_fd_sc_hd__or2_4
XFILLER_0_8_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_115_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08223_ _04094_ _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09588__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _04005_ _04038_ _04037_ _04009_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08796__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08085_ _03947_ net225 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1136_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12380__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09760__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net883 _04639_ _04651_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] _03816_ net262 vssd1 vssd1
+ vccd1 vccd1 _03829_ sky130_fd_sc_hd__or3b_1
X_16765__1319 vssd1 vssd1 vccd1 vccd1 _16765__1319/HI net1319 sky130_fd_sc_hd__conb_1
XANTENNA__10107__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09512__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07869_ _03758_ _03759_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__or2_2
XANTENNA__15597__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11724__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[16\] net688 net664 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10880_ net382 _06071_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] net721 net710 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a221o_1
XANTENNA__13224__B net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12550_ net286 net2139 net466 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11501_ net418 _06743_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ net319 net2118 net482 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__mux2_1
XANTENNA__12555__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ net1018 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XANTENNA__09579__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _06098_ _06102_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ net1152 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XANTENNA__16222__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ net459 team_02_WB.instance_to_wrap.top.aluOut\[11\] _06974_ _06887_ vssd1
+ vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__o22a_4
XANTENNA__10594__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13102_ net230 _03109_ net228 _07091_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_131_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] net724 net720 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a22o_1
X_14082_ net1091 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
X_11294_ net461 team_02_WB.instance_to_wrap.top.aluOut\[14\] _06911_ _06887_ vssd1
+ vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__o22a_4
X_13033_ _03050_ _03051_ _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12290__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ _05896_ _05897_ _05899_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_1512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11543__C1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1104 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1111 net1113 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
XANTENNA__09165__A _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1122 net1137 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
X_10176_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] net732 net720 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__a22o_1
XANTENNA__09751__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1133 net1137 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_2
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_4
Xfanout1155 net1160 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__buf_2
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_4
X_14984_ net1047 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__C1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1177 net1180 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
Xfanout1188 net1189 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1199 net1202 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_2
XANTENNA__09503__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16723_ net1277 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
X_13935_ net1127 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16654_ net1388 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ net1050 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672__1227 vssd1 vssd1 vccd1 vccd1 _16672__1227/HI net1227 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15605_ clknet_leaf_115_wb_clk_i _02056_ _00563_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12817_ _07391_ _07440_ _07392_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16585_ clknet_leaf_81_wb_clk_i net1408 _01458_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13797_ net1073 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15536_ clknet_leaf_41_wb_clk_i _01987_ _00494_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12748_ _04846_ _06231_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12810__A2 _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10821__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15467_ clknet_leaf_20_wb_clk_i _01918_ _00425_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12679_ _07292_ _07295_ _07298_ _07306_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__or4b_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14418_ net1085 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15398_ clknet_leaf_12_wb_clk_i _01849_ _00356_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11377__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14349_ net1134 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09059__B _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold638 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09990__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08910_ net973 _04407_ _03396_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__mux2_1
XANTENNA__11809__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16019_ clknet_leaf_125_wb_clk_i _02470_ _00977_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09890_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\] net763 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\]
+ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a221o_1
XANTENNA__10337__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ net15 net949 net923 net2379 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XANTENNA__10888__A1 _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1305 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[6\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[6\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__mux2_2
Xhold1338 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 team_02_WB.instance_to_wrap.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net2747
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07723_ _03612_ _03613_ _03611_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07654_ _03509_ _03537_ _03513_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09522__B _05193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08419__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07585_ _03474_ _03475_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout344_A _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1086_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[23\] net666 net655 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a22o_1
XANTENNA__11065__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12793__A_N _05797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09255_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] net808 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[25\]
+ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12375__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout511_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ _04035_ _04039_ _04059_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__mux2_4
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09186_ net898 _04865_ _04630_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a21o_1
XANTENNA__08769__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ _04017_ _04019_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10040__A2 _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08068_ _03900_ _03935_ _03936_ _03897_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09981__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16521__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\] net809 net801 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a22o_1
XANTENNA__09194__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16740__1294 vssd1 vssd1 vccd1 vccd1 _16740__1294/HI net1294 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ net2171 net296 net532 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13720_ net1056 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
X_10932_ net391 _06406_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__or2_1
XANTENNA__08329__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ net1127 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
X_10863_ _06411_ _06509_ net450 vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__o21a_1
X_12602_ _07019_ _07050_ _07059_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__or4_1
X_16370_ clknet_leaf_74_wb_clk_i _00011_ _01262_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.noisy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11056__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13582_ net1150 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10794_ _06060_ _06070_ net376 vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12793__B _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15321_ clknet_leaf_106_wb_clk_i _01772_ _00279_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12533_ net238 net2630 net466 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12285__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ clknet_leaf_52_wb_clk_i _01703_ _00210_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15612__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ net361 net2246 net484 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14203_ net1047 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _06941_ _07021_ net386 vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__mux2_1
X_15183_ clknet_leaf_34_wb_clk_i _01634_ _00141_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12395_ net345 net2424 net494 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__mux2_1
XANTENNA__10567__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ net1106 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XANTENNA__10031__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _06091_ _06094_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11629__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ net1029 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
X_11277_ _06847_ _06895_ net380 vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__mux2_1
XANTENNA__10319__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ team_02_WB.instance_to_wrap.top.pc\[20\] net944 net941 _03038_ vssd1 vssd1
+ vccd1 vccd1 _01518_ sky130_fd_sc_hd__a22o_1
X_10228_ net398 _05882_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__nor2_1
XANTENNA__09724__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08932__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[18\] vssd1 vssd1 vccd1 vccd1
+ net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net897 _05797_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o21a_1
XANTENNA__16118__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ net1034 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XANTENNA__10769__A _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ net1260 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13918_ net1070 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14898_ net1147 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13849_ net1060 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_16637_ net1208 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XANTENNA__15142__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16568_ clknet_leaf_99_wb_clk_i net1423 _01441_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08999__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15519_ clknet_leaf_24_wb_clk_i _01970_ _00477_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12195__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16499_ clknet_leaf_0_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[2\]
+ _01373_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15292__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net854 net770 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10270__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16764__1318 vssd1 vssd1 vccd1 vccd1 _16764__1318/HI net1318 sky130_fd_sc_hd__conb_1
XFILLER_0_83_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold402 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold413 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10022__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold424 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08620__C1 _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold435 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold468 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ _05598_ _05600_ _05602_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold479 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_2
Xfanout926 net927 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09715__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\] net690 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\]
+ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a221o_1
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_2
Xfanout948 _04554_ vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A _06935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 _04273_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__buf_2
X_08824_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net6 vssd1 vssd1 vccd1 vccd1
+ _04554_ sky130_fd_sc_hd__nand2_1
Xhold1102 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 net109 vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1135 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net1619 net956 net925 _04534_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
Xhold1157 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout461_A _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1179 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout559_A _07197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _03551_ _03591_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ net748 _04446_ _04466_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07637_ _03494_ _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or2_1
XANTENNA__13027__A2 _07336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout726_A _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07568_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03457_ team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15635__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold137_A team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] net794 _04975_ _04984_
+ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16516__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] net2746 net969 vssd1
+ vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09238_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[25\] net697 net665 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\]
+ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a221o_1
XANTENNA__10261__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\] net866 net774 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ net455 _06185_ _06821_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11210__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net297 net2244 net516 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
XANTENNA__09954__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16671__1226 vssd1 vssd1 vccd1 vccd1 _16671__1226/HI net1226 sky130_fd_sc_hd__conb_1
XFILLER_0_82_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _06058_ _06069_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold980 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09167__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09706__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _06340_ _06695_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] net736 net704 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ clknet_leaf_12_wb_clk_i _02321_ _00828_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08758__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A wbm_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1199 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14752_ net1182 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11964_ net353 net2015 net536 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ net1134 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
X_10915_ _06239_ _06306_ _06236_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14683_ net1194 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_11895_ net349 net2351 net546 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XANTENNA__08693__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output109_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11912__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16422_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[21\]
+ _01296_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_13634_ net1090 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
X_10846_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16560__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ clknet_leaf_102_wb_clk_i _02786_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13565_ net1173 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__inv_2
XANTENNA__13412__B _03297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777_ net415 net436 _06418_ net453 _04744_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a32o_1
XANTENNA__10788__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15304_ clknet_leaf_86_wb_clk_i _01755_ _00262_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12516_ net2012 net268 net476 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ clknet_leaf_101_wb_clk_i _02717_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13496_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] _03176_ _03345_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15235_ clknet_leaf_43_wb_clk_i _01686_ _00193_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12447_ net315 net2167 net485 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10004__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09945__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15166_ clknet_leaf_3_wb_clk_i _01617_ _00124_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12378_ net287 net2488 net492 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14117_ net1087 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11329_ net402 _06942_ _06943_ net409 vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__o211a_1
X_15097_ clknet_leaf_112_wb_clk_i _01548_ _00055_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09158__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14048_ net1083 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15999_ clknet_leaf_27_wb_clk_i _02450_ _00957_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_08540_ net84 net2698 net893 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ _03420_ _04284_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09881__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__B2 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10243__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09023_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\] net688 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\]
+ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout307_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 net138 vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 net126 vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold232 team_02_WB.instance_to_wrap.top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1 net1630
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold243 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold265 team_02_WB.START_ADDR_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_02_WB.instance_to_wrap.top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1
+ net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold287 team_02_WB.instance_to_wrap.top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1 net1685
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 net703 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09149__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09925_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] net734 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a22o_1
Xfanout712 _04457_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_6
Xhold298 team_02_WB.instance_to_wrap.top.pc\[12\] vssd1 vssd1 vccd1 vccd1 net1696
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout723 _04453_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_2
XANTENNA__15188__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 _04447_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_6
Xfanout745 _04441_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 _04680_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_4
X_09856_ _05508_ _05516_ _05518_ _05520_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[11\]
+ sky130_fd_sc_hd__or4_4
Xfanout767 _04674_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
Xfanout778 _04670_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
XANTENNA__07482__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 net792 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
X_08807_ net157 net952 net903 net1533 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
X_09787_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[12\] net738 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\]
+ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout843_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08738_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[23\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[23\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09321__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08675__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11732__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ _05052_ net367 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nand2_1
XANTENNA__12208__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net295 net2339 net568 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
XANTENNA__08607__A team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _06269_ _06281_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16824__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10234__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ team_02_WB.instance_to_wrap.top.a1.row1\[18\] _03222_ _03240_ team_02_WB.instance_to_wrap.top.a1.row2\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a22o_1
X_10562_ _04723_ _04741_ _06214_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ _04576_ _07190_ _07194_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__or3_4
XFILLER_0_107_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13281_ _03182_ _03185_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__nor2_1
XANTENNA__12563__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _05614_ _06016_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15020_ net1190 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
X_12232_ net352 net2548 net512 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__mux2_1
XANTENNA__09438__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net342 net2389 net520 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ _05156_ net453 net451 _06744_ _06742_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ net336 net1905 net524 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11907__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _06564_ _06679_ net384 vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__mux2_1
X_15922_ clknet_leaf_10_wb_clk_i _02373_ _00880_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09560__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15800__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ clknet_leaf_21_wb_clk_i _02304_ _00811_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_16763__1317 vssd1 vssd1 vccd1 vccd1 _16763__1317/HI net1317 sky130_fd_sc_hd__conb_1
X_14804_ net1199 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15784_ clknet_leaf_85_wb_clk_i _02235_ _00742_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12996_ _07451_ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12998__A1 team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14735_ net1040 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
X_11947_ net304 net2363 net538 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15950__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14666_ net1041 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ net280 net2143 net544 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16405_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[4\]
+ _01279_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] sky130_fd_sc_hd__dfrtp_4
X_13617_ net1030 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
X_10829_ net911 _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14597_ net1198 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11422__A1 _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ _03383_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16336_ clknet_leaf_100_wb_clk_i _02769_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09091__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16267_ clknet_leaf_93_wb_clk_i _02700_ _01219_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12473__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03132_ vssd1 vssd1 vccd1
+ vccd1 _03342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09379__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ clknet_leaf_21_wb_clk_i _01669_ _00176_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16198_ clknet_leaf_96_wb_clk_i _02643_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15149_ clknet_leaf_32_wb_clk_i _01600_ _00107_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07971_ _03831_ _03834_ _03858_ _03859_ _03839_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11817__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ _05368_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__nor2_8
XANTENNA__11489__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15480__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\] net769 _05308_ _05310_
+ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net695 net687 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09303__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ net63 net62 net59 net60 vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout257_A _06553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16670__1225 vssd1 vssd1 vccd1 vccd1 _16670__1225/HI net1225 sky130_fd_sc_hd__conb_1
X_08454_ _04310_ net1651 _04286_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08385_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] _04254_ _04255_ vssd1 vssd1
+ vccd1 vccd1 _04257_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12891__B _05797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] net793 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout793_A _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09790__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15823__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout520 _07212_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout531 _07209_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11727__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 _07202_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09908_ _05543_ _05569_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__and2_1
Xfanout553 net555 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout564 _07195_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_6
Xfanout575 _07191_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_4
Xfanout586 _07211_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09839_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[11\] net800 net784 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a22o_1
XANTENNA__13227__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ team_02_WB.instance_to_wrap.top.pc\[26\] _06238_ vssd1 vssd1 vccd1 vccd1
+ _02884_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _07192_ _07194_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12558__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05678_ _05681_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__and2_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14339__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14520_ net1105 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11732_ net351 net2146 net564 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
XANTENNA__15203__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14451_ net1128 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
X_11663_ net356 net2403 net575 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ net1479 _04267_ net828 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
X_10614_ net750 _05795_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__o21a_2
XANTENNA__10207__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ net1114 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09073__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ _07183_ _07184_ _07171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[0\]
+ sky130_fd_sc_hd__nand3b_2
XFILLER_0_84_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16121_ clknet_leaf_64_wb_clk_i _02567_ _01079_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ _03218_ _03231_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__nor2_2
XFILLER_0_52_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12293__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _06197_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ clknet_leaf_51_wb_clk_i _02503_ _01010_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ _03175_ _03176_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[11\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__a211o_1
X_10476_ _04603_ _06128_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nor2_1
X_15003_ net1166 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12215_ net306 net2205 net515 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ team_02_WB.START_ADDR_VAL_REG\[3\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net217 sky130_fd_sc_hd__a21o_1
XFILLER_0_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14802__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09781__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net287 net2333 net520 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11637__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12077_ net277 net2372 net525 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15905_ clknet_leaf_5_wb_clk_i _02356_ _00863_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11028_ _05053_ _05072_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15836_ clknet_leaf_50_wb_clk_i _02287_ _00794_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12468__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ _07454_ _03005_ net888 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15767_ clknet_leaf_119_wb_clk_i _02218_ _00725_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14718_ net1033 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15698_ clknet_leaf_15_wb_clk_i _02149_ _00656_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14649_ net1003 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08170_ _04023_ _04032_ _04020_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09064__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16319_ clknet_leaf_96_wb_clk_i _02752_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08811__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__10017__A _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 wbm_stb_o sky130_fd_sc_hd__buf_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07954_ _03805_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07885_ _03706_ _03736_ _03707_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__o21a_1
XANTENNA__10134__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\] net704 net701 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a221o_1
XANTENNA__15226__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _05220_ _05222_ _05224_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12378__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A _07202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08506_ _04279_ _04325_ _04336_ _04337_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[19\] net711 net666 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a22o_1
XANTENNA__15376__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ net960 _04285_ _04297_ _04298_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16621__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08368_ _04232_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nand2_2
XFILLER_0_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08802__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08299_ _04161_ _04166_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__xor2_2
XANTENNA__10070__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16762__1316 vssd1 vssd1 vccd1 vccd1 _16762__1316/HI net1316 sky130_fd_sc_hd__conb_1
XFILLER_0_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[0\] net877 net772 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10261_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\] net688 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12000_ net1845 net360 net532 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
X_10192_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\] net808 net792 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\]
+ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a221o_1
XANTENNA__16001__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout350 _03645_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout361 _07170_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09515__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_2
X_13951_ net1125 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
Xfanout383 net385 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
Xfanout394 net397 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _02926_ _02935_ _02924_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o21a_1
X_13882_ net1045 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
X_16670_ net1225 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__16151__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08766__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12796__B _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ _04889_ _06235_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a21o_1
X_15621_ clknet_leaf_125_wb_clk_i _02072_ _00579_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12288__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12764_ _05247_ _05256_ _06260_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__or3_1
X_15552_ clknet_leaf_9_wb_clk_i _02003_ _00510_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14503_ net1136 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
X_11715_ net306 net2155 net567 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15483_ clknet_leaf_104_wb_clk_i _01934_ _00441_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12695_ _04435_ _04592_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__nor2_1
XANTENNA__11920__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11646_ net295 net1989 net572 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
X_14434_ net1093 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09046__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15869__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 wbm_dat_i[16] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput25 wbm_dat_i[26] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1055 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
Xinput36 wbm_dat_i[7] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] net887 _07168_ team_02_WB.instance_to_wrap.top.pc\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput47 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_16104_ clknet_leaf_70_wb_clk_i _02550_ _01062_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13316_ net987 _03221_ net986 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__and3b_1
Xinput69 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10521__A_N _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10528_ _06149_ _06178_ _06180_ _06150_ _06177_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__o221a_1
X_14296_ net1063 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
Xhold809 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16035_ clknet_leaf_45_wb_clk_i _02486_ _00993_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13247_ net1664 net980 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10459_ _04502_ net374 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _03150_ _03153_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__nor2_1
X_12129_ net346 net2127 net588 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09506__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07670_ _03531_ _03556_ _03524_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__and3b_1
XANTENNA_wire607_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15819_ clknet_leaf_19_wb_clk_i _02270_ _00777_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15399__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ net1353 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
X_09340_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[23\] net820 net848 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10300__A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ _04943_ _04945_ _04947_ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__or4_1
X_16709__1263 vssd1 vssd1 vccd1 vccd1 _16709__1263/HI net1263 sky130_fd_sc_hd__conb_1
XFILLER_0_34_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11830__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14707__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _04079_ _04093_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ _04008_ _04036_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08424__B net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08084_ _03941_ _03969_ _03970_ _03937_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__o22a_2
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16024__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1129_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__B1 _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08986_ net883 _04636_ _04644_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__and3_2
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07937_ _03409_ net262 _03816_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07868_ _03732_ _03757_ _03723_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07490__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07799_ _03675_ _03689_ net341 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__o21a_1
X_09538_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[18\] net737 net645 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09276__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\] net874 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08484__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11740__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11500_ net394 _06942_ _07098_ net411 vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__o211a_1
XANTENNA__10291__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12480_ net315 net2265 net481 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__mux2_1
XANTENNA__10830__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10544__A_N _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13240__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ _05703_ _06166_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14150_ net1092 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ team_02_WB.instance_to_wrap.top.pc\[11\] net908 _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[11\]
+ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ _02926_ _02935_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] net692 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\]
+ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14081_ net1144 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XANTENNA__12571__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11293_ _06268_ net743 _06909_ _06281_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13032_ net231 _03049_ net228 _06828_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09736__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] net869 net793 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\]
+ _05894_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__a221o_1
XANTENNA__09200__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1101 net1104 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_2
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] net657 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\]
+ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a221o_1
XANTENNA__10897__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1123 net1126 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net1136 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_2
Xfanout1156 net1159 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
X_14983_ net1035 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15541__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1180 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
XANTENNA__11915__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1192 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_2
X_16722_ net1276 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
X_13934_ net1116 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12600__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ net1220 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_13865_ net1011 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15604_ clknet_leaf_51_wb_clk_i _02055_ _00562_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12816_ _05379_ _06268_ _07439_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__a21o_1
X_16584_ clknet_leaf_85_wb_clk_i net1406 _01457_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09267__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13796_ net1101 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ clknet_leaf_32_wb_clk_i _01986_ _00493_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _04846_ _06231_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11650__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10282__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15466_ clknet_leaf_46_wb_clk_i _01917_ _00424_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12678_ _06920_ _06945_ _07299_ _07305_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11629_ net356 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\] net579 vssd1
+ vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XANTENNA__13150__B _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14417_ net1078 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
XANTENNA__13220__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15397_ clknet_leaf_127_wb_clk_i _01848_ _00355_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10034__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09975__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ net1004 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold606 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold617 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14279_ net1153 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XANTENNA__12481__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09727__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09356__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ clknet_leaf_10_wb_clk_i _02469_ _00976_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08840_ net16 net949 net923 team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1
+ vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XANTENNA__10888__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1306 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ net1584 net958 net926 _04542_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
Xhold1317 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1328 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11825__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _03582_ _03606_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__xor2_2
XFILLER_0_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13606__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16761__1315 vssd1 vssd1 vccd1 vccd1 _16761__1315/HI net1315 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07584_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] _03470_ _03471_ vssd1 vssd1
+ vccd1 vccd1 _03475_ sky130_fd_sc_hd__and3_1
XANTENNA__09258__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09323_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[23\] net727 net694 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11560__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\] net779 net768 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1079_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08205_ _04083_ _04087_ _04064_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a21o_2
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13211__B1 _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ _04865_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[27\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout504_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10025__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__B2 _04541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _04013_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__or2_1
XANTENNA__09966__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09430__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08067_ _03922_ _03953_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12391__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07485__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09718__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15564__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ _04653_ net886 _04637_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ net2225 net287 net532 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09497__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10931_ _06395_ _06402_ net391 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__mux2_1
XANTENNA__13235__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10862_ net420 _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__nor2_1
X_13650_ net1081 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09249__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12601_ _07078_ _07104_ _07228_ _07128_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__or4b_1
XFILLER_0_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11056__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13581_ net1170 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12566__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ net363 _06065_ _06066_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12532_ net594 _07207_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__nand2_4
XFILLER_0_82_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10264__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15320_ clknet_leaf_124_wb_clk_i _01771_ _00278_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08899__B1_N net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12463_ net353 net2334 net484 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
X_15251_ clknet_leaf_3_wb_clk_i _01702_ _00209_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13202__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202_ net1038 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_11414_ _06979_ _07020_ net380 vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__mux2_1
XANTENNA__09957__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15182_ clknet_leaf_40_wb_clk_i _01633_ _00140_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12394_ net347 net1780 net494 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09421__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ net1119 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XANTENNA__12961__C1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _06019_ _06148_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14082__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14064_ net1021 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11276_ _06360_ _06383_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ _06748_ net226 _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10227_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__inv_2
X_16708__1262 vssd1 vssd1 vccd1 vccd1 _16708__1262/HI net1262 sky130_fd_sc_hd__conb_1
XANTENNA__09904__A _05567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[4\] vssd1 vssd1 vccd1
+ vccd1 _05815_ sky130_fd_sc_hd__or2_1
Xhold3 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[13\] vssd1 vssd1 vccd1 vccd1
+ net1401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11645__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ _05722_ _05745_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__and2_1
X_14966_ net1010 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09488__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ net1259 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_37_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ net1105 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14897_ net1171 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ net1207 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_13848_ net1107 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16567_ clknet_leaf_99_wb_clk_i net1427 _01440_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12476__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13779_ net1148 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10255__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15518_ clknet_leaf_3_wb_clk_i _01969_ _00476_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16498_ clknet_leaf_7_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[1\]
+ _01372_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09660__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15449_ clknet_leaf_106_wb_clk_i _01900_ _00407_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10007__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09412__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15587__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold403 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold414 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold436 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold447 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09941_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] net871 net795 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[9\]
+ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a221o_1
Xhold469 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_2
Xfanout916 _04278_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_2
Xfanout927 _04517_ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
X_09872_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\] net666 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a22o_1
Xfanout938 _03422_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_2
Xfanout949 _04553_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
X_08823_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net6 vssd1 vssd1 vccd1 vccd1
+ _04553_ sky130_fd_sc_hd__and2_1
Xhold1103 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1136 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[15\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[15\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__mux2_1
Xhold1158 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07705_ _03586_ _03589_ _03593_ _03594_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08685_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] net660 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07636_ _03489_ _03491_ _03492_ _03506_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__or4b_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12894__B _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07567_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] team_02_WB.instance_to_wrap.top.a1.dataIn\[28\]
+ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__or3_1
XANTENNA__11038__A2 team_02_WB.instance_to_wrap.top.aluOut\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12386__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A _04495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09306_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net854 net802 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a22o_1
XANTENNA__10246__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09100__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07498_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] team_02_WB.instance_to_wrap.ramload\[7\]
+ net967 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16362__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09651__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09237_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[25\] net638 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09939__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\] net863 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ _03999_ _04002_ _04004_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__A2 team_02_WB.instance_to_wrap.top.aluOut\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09099_ _04768_ _04769_ _04778_ _04781_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[29\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_124_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _06757_ _06758_ net411 vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold981 team_02_WB.instance_to_wrap.ramload\[17\] vssd1 vssd1 vccd1 vccd1 net2379
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold992 team_02_WB.instance_to_wrap.top.pad.keyCode\[1\] vssd1 vssd1 vccd1 vccd1
+ net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ team_02_WB.instance_to_wrap.top.pc\[21\] _06339_ team_02_WB.instance_to_wrap.top.pc\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\] net693 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\]
+ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13246__A team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14820_ net1202 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08390__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input15_A wbm_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14751_ net1182 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
X_11963_ net356 net1951 net538 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13702_ net1092 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ _06235_ _06323_ net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] net443
+ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a221o_1
X_14682_ net1167 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
X_11894_ net338 net2549 net546 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XANTENNA__08774__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09890__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16421_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[20\]
+ _01295_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10845_ net365 _06405_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__nor2_1
X_13633_ net1101 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XANTENNA__12296__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10237__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16352_ clknet_leaf_96_wb_clk_i _02785_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10776_ _06414_ _06423_ net450 vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__o21a_1
X_13564_ net1173 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__inv_2
XANTENNA__10788__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09642__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15303_ clknet_leaf_15_wb_clk_i _01754_ _00261_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ net1697 net323 net476 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08850__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13495_ net2165 _03350_ _03351_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__o21a_1
X_16283_ clknet_leaf_101_wb_clk_i _02716_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ clknet_leaf_50_wb_clk_i _01685_ _00192_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12446_ net303 net2310 net487 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ clknet_leaf_113_wb_clk_i _01616_ _00123_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12377_ net279 net2581 net492 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__mux2_1
X_16760__1314 vssd1 vssd1 vccd1 vccd1 _16760__1314/HI net1314 sky130_fd_sc_hd__conb_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11328_ net395 _06737_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__or2_1
X_14116_ net1093 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15096_ clknet_leaf_121_wb_clk_i _01547_ _00054_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14047_ net1121 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
X_11259_ net418 _06117_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12783__A_N _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15998_ clknet_leaf_3_wb_clk_i _02449_ _00956_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14949_ net1047 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08470_ _04322_ net1698 net827 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ clknet_leaf_62_wb_clk_i _02853_ _01492_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09094__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10779__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09633__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\] net733 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08652__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 net122 vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold211 _02637_ vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 net177 vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08432__B net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 team_02_WB.START_ADDR_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold244 team_02_WB.START_ADDR_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_02_WB.instance_to_wrap.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net1664
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_02_WB.instance_to_wrap.top.a1.row1\[109\] vssd1 vssd1 vccd1 vccd1 net1675
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_02_WB.instance_to_wrap.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net1686
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold299 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\] net682 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a221o_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_6
Xfanout713 _04457_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1111_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 _04450_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_6
Xfanout735 _04447_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_2
Xfanout746 _04441_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09544__A _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A wbm_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[11\] net776 net844 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout757 _04679_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout571_A _07193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _04674_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_4
Xfanout779 _04670_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout669_A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net158 net952 net904 net1536 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
X_09786_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\] net718 net702 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08737_ net1662 net955 net924 _04525_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout836_A _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08668_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\] net705 _04464_ vssd1
+ vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09872__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ _03406_ _03506_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__xnor2_2
XANTENNA__16527__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _04380_ _04393_ _04386_ _04376_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15752__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__B net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16664__1398 vssd1 vssd1 vccd1 vccd1 net1398 _16664__1398/LO sky130_fd_sc_hd__conb_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10630_ team_02_WB.instance_to_wrap.top.pc\[15\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _06282_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09085__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09624__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11967__B1 _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16707__1261 vssd1 vssd1 vccd1 vccd1 _16707__1261/HI net1261 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _04744_ _06213_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__nor2_1
XANTENNA__08832__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net235 net2355 net505 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _03179_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10492_ _05075_ _06040_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ net354 net1955 net515 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ net346 net1834 net521 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11113_ net416 _06743_ _06412_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__o21ai_1
X_12093_ net331 net2433 net526 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12799__B _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ _06631_ _06678_ net379 vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__mux2_1
X_15921_ clknet_leaf_18_wb_clk_i _02372_ _00879_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15852_ clknet_leaf_22_wb_clk_i _02303_ _00810_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07571__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10170__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ net1201 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ clknet_leaf_15_wb_clk_i _02234_ _00741_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12995_ _07377_ _07378_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__nand2_1
XANTENNA__11923__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14734_ net1040 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12998__A2 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11946_ net298 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] net536 vssd1
+ vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09863__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14665_ net1043 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ net273 net2323 net546 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16404_ clknet_leaf_75_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[3\]
+ _01278_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_131_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13616_ net1003 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XANTENNA__09076__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10828_ team_02_WB.instance_to_wrap.top.pc\[29\] _06344_ vssd1 vssd1 vccd1 vccd1
+ _06476_ sky130_fd_sc_hd__xnor2_1
X_14596_ net1198 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XANTENNA__09615__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16335_ clknet_leaf_100_wb_clk_i _02768_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_13547_ _03385_ _03386_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14535__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10759_ net408 _06365_ _06381_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16266_ clknet_leaf_96_wb_clk_i _00004_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_13478_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\] _03132_ vssd1 vssd1 vccd1
+ vccd1 _03341_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15217_ clknet_leaf_17_wb_clk_i _01668_ _00175_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12429_ net355 net2472 net491 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__mux2_1
X_16197_ clknet_leaf_70_wb_clk_i net1498 _01155_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ clknet_leaf_23_wb_clk_i _01599_ _00106_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07970_ net2675 net936 net919 _03860_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a22o_1
X_15079_ clknet_leaf_80_wb_clk_i _01530_ _00042_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15625__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09000__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09640_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[16\] net777 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\]
+ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10161__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[17\] net739 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\]
+ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08522_ net46 net49 net48 net47 vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or4b_1
XFILLER_0_37_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11833__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09854__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ net960 _04308_ _04309_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13399__C1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08384_ _04254_ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08814__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1061_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09005_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\] net817 net849 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout786_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout510 _07216_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_6
XFILLER_0_121_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09274__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 _07212_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
X_09907_ _05543_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout532 net535 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_6
Xfanout543 _07202_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout565 _07195_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_4
Xfanout576 net579 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout587 _07211_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_4
X_09838_ _05493_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__nor2_4
XFILLER_0_96_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07553__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09769_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] net761 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11743__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11800_ net233 net2345 net559 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__and2b_1
XANTENNA__09845__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11731_ net357 net1874 net567 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
XANTENNA__13243__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14450_ net1082 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11662_ net342 net2490 net572 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13401_ net1484 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] _03297_ vssd1 vssd1
+ vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10613_ net929 _05841_ _06220_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a21o_1
X_14381_ net1133 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XANTENNA__12574__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _04598_ _04602_ _04702_ _06217_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__or4_1
X_16120_ clknet_leaf_62_wb_clk_i _02566_ _01078_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input82_A wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ _05094_ _05113_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2b_1
X_13332_ net987 _03208_ net986 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__and3b_1
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16080__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16051_ clknet_leaf_126_wb_clk_i _02502_ _01009_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13263_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[8\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _03176_
+ sky130_fd_sc_hd__and3_1
X_10475_ _04584_ _04596_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15002_ net1189 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XANTENNA__15648__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12214_ net295 net2452 net512 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__mux2_1
X_13194_ team_02_WB.START_ADDR_VAL_REG\[2\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net214 sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ net279 net2163 net520 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
XANTENNA__11918__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07792__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12076_ net263 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[25\] net526 vssd1
+ vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux2_1
X_11027_ _05075_ _06663_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__nor2_1
X_15904_ clknet_leaf_11_wb_clk_i _02355_ _00862_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10143__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15835_ clknet_leaf_104_wb_clk_i _02286_ _00793_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11653__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09297__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15766_ clknet_leaf_86_wb_clk_i _02217_ _00724_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12978_ _07454_ _03005_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__or2_1
XANTENNA__09836__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14717_ net1035 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11929_ net344 net2152 net541 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
X_15697_ clknet_leaf_16_wb_clk_i _02148_ _00655_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09049__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14648_ net1001 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15178__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12484__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16423__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14579_ net1145 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10603__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16318_ clknet_leaf_97_wb_clk_i _02751_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16249_ clknet_leaf_93_wb_clk_i _02687_ _01206_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[13] sky130_fd_sc_hd__buf_2
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[23] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__11828__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16663__1397 vssd1 vssd1 vccd1 vccd1 net1397 _16663__1397/LO sky130_fd_sc_hd__conb_1
X_07953_ _03824_ net262 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nand2_1
X_16706__1260 vssd1 vssd1 vccd1 vccd1 _16706__1260/HI net1260 sky130_fd_sc_hd__conb_1
X_07884_ _03751_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__or3_1
XANTENNA__10134__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07535__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[16\] net676 net672 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\] net834 net754 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[18\]
+ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__a221o_1
XANTENNA__09288__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09827__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__B2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11095__B1 team_02_WB.instance_to_wrap.top.aluOut\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _04325_ team_02_WB.instance_to_wrap.top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1
+ _04337_ sky130_fd_sc_hd__and2b_1
X_09485_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\] net702 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout534_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ net2723 _04286_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08367_ _03410_ _04228_ _04221_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12394__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout701_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07488__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _04166_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__or2_2
XFILLER_0_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08015__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10260_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] net668 _05914_ vssd1
+ vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a21o_1
XANTENNA__09212__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\] net800 net836 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11570__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__B2 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout340 _07075_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_2
Xfanout351 _07153_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_2
Xfanout362 _03568_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13950_ net1022 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
Xfanout373 net375 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_2
XANTENNA__10125__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net397 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlymetal6s2s_1
X_12901_ team_02_WB.instance_to_wrap.top.pc\[4\] _05843_ _02934_ vssd1 vssd1 vccd1
+ vccd1 _02935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09732__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ net1058 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XANTENNA__12569__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15620_ clknet_leaf_54_wb_clk_i _02071_ _00578_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12832_ _07374_ _02865_ _07373_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09279__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13075__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13075__B2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15551_ clknet_leaf_27_wb_clk_i _02002_ _00509_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12763_ _05215_ _06257_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15320__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14502_ net1139 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11714_ net295 net2434 net564 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XANTENNA__08782__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15482_ clknet_leaf_119_wb_clk_i _01933_ _00440_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12694_ _07238_ _07251_ _07321_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__and3_1
X_14433_ net1102 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
X_11645_ net289 net2682 net572 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
XANTENNA__12586__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15470__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput15 wbm_dat_i[17] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14364_ net1123 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
Xinput26 wbm_dat_i[27] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ _04581_ _06325_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__and2b_1
XANTENNA__09451__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput37 wbm_dat_i[8] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_2
XFILLER_0_68_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput48 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_16103_ clknet_leaf_71_wb_clk_i _02549_ _01061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput59 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ _03214_ _03397_ team_02_WB.instance_to_wrap.top.lcd.nextState\[4\] vssd1
+ vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__and3b_2
X_10527_ _05572_ _06147_ _06174_ _06179_ _06172_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__o311a_1
X_14295_ net1108 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XANTENNA__14813__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16034_ clknet_leaf_50_wb_clk_i _02485_ _00992_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ team_02_WB.instance_to_wrap.ramload\[19\] net980 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[19\] sky130_fd_sc_hd__and2_1
X_10458_ _05975_ net370 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and2_1
XANTENNA__09907__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11648__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ _03161_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__nor2_1
X_10389_ _04993_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12128_ net339 net1941 net588 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12059_ net327 net2068 net530 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10116__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12479__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13164__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ clknet_leaf_44_wb_clk_i _02269_ _00776_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ net1352 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
XANTENNA__09809__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15749_ clknet_leaf_127_wb_clk_i _02200_ _00707_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10300__B team_02_WB.instance_to_wrap.top.DUT.read_data2\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] net863 net786 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\]
+ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _04076_ _04092_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08152_ _04025_ _04032_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09442__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08083_ _03939_ _03950_ net225 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08796__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15963__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09817__A _05461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _04640_ _04653_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout484_A _07222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ _03409_ net262 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10107__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07867_ _03723_ _03732_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__and3_2
XANTENNA__12389__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16469__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__A2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ _05257_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07798_ _03676_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__and2_1
XANTENNA__13057__B2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09537_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\] net633 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[18\]
+ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\] net841 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a22o_1
XANTENNA__09681__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08419_ net919 _04268_ _04283_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or3_2
XFILLER_0_136_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09399_ _05052_ _05072_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11430_ net332 net1892 net584 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09433__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11361_ net913 _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ _07408_ _07419_ _07421_ net890 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__o31ai_1
X_10312_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\] net712 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14080_ net1075 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
X_11292_ net913 _06908_ _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1
+ vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_132_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08631__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _07388_ _07389_ _07443_ net888 vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a31o_1
X_10243_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[2\] net809 net805 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\]
+ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a221o_1
XANTENNA_input45_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] net712 net670 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a22o_1
Xfanout1102 net1104 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1113 net1137 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_2
XFILLER_0_100_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1124 net1126 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
Xfanout1135 net1136 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_4
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_2
Xfanout1157 net1159 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_2
X_14982_ net1044 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__A1 team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__buf_4
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_2
X_16721_ net1275 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
X_13933_ net1133 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XANTENNA__12299__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ net1219 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13864_ net1100 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ clknet_leaf_3_wb_clk_i _02054_ _00561_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ _07393_ _07394_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16583_ clknet_leaf_87_wb_clk_i net1410 _01456_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ net1075 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11931__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14808__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15534_ clknet_leaf_42_wb_clk_i _01985_ _00492_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _04804_ _06228_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09672__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15465_ clknet_leaf_29_wb_clk_i _01916_ _00423_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_16662__1396 vssd1 vssd1 vccd1 vccd1 net1396 _16662__1396/LO sky130_fd_sc_hd__conb_1
X_12677_ _06878_ _07301_ _07302_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__and4_1
X_14416_ net1006 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11628_ net344 net2635 net577 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15396_ clknet_leaf_55_wb_clk_i _01847_ _00354_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09424__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14347_ net1025 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[2\] _07152_ vssd1 vssd1 vccd1
+ vccd1 _07153_ sky130_fd_sc_hd__a21o_4
XFILLER_0_53_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15216__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold618 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ net1142 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16017_ clknet_leaf_111_wb_clk_i _02468_ _00975_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13229_ team_02_WB.instance_to_wrap.ramload\[2\] net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_42_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10337__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1307 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16611__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1318 team_02_WB.instance_to_wrap.top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 net2716
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[7\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[7\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1329 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
X_07721_ team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] _03606_ _03607_ vssd1 vssd1
+ vccd1 vccd1 _03612_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ _03510_ _03539_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13039__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ _03470_ _03471_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1
+ vccd1 vccd1 _03474_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11841__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] net714 net675 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09663__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09253_ _04922_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ _04083_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ _04855_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09415__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ _03981_ _04012_ _03978_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _03923_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10328__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout866_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__B team_02_WB.instance_to_wrap.top.DUT.read_data2\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] net886 net882 _04635_
+ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ _03789_ _03792_ _03767_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o21a_1
XANTENNA__11421__A2_N _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08899_ _04398_ _04408_ net910 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ net399 _06570_ _06571_ _06572_ net416 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_92_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10861_ _06413_ _06420_ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11751__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net440 _07160_ _07178_ _07144_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ net1150 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08626__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ net363 _06083_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nor2_1
XANTENNA__09654__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12531_ net1800 net235 net477 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15239__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15250_ clknet_leaf_10_wb_clk_i _01701_ _00208_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12462_ net354 net2364 net487 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14201_ net1061 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11413_ _06389_ _06392_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__nand2_1
X_15181_ clknet_leaf_23_wb_clk_i _01632_ _00139_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12582__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12393_ net337 net1859 net494 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14132_ net1037 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11344_ _06147_ _06860_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ net1129 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
X_11275_ _06025_ _06893_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10319__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ net232 _03036_ _07448_ _03034_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10226_ _05872_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__nor2_4
XFILLER_0_20_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08393__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _05801_ _05810_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[4\]
+ sky130_fd_sc_hd__or4_4
Xhold4 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[29\] vssd1 vssd1 vccd1 vccd1
+ net1402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14965_ net1002 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
X_10088_ _05722_ _05745_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16704_ net1258 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
X_13916_ net1124 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14896_ net1172 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16635_ net1383 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XANTENNA__16014__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13847_ net1112 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11661__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16566_ clknet_leaf_81_wb_clk_i net1447 _01439_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13778_ net1078 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08999__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15517_ clknet_leaf_111_wb_clk_i _01968_ _00475_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12729_ net961 _04279_ _03418_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16497_ clknet_leaf_6_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[0\]
+ _01371_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16164__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15448_ clknet_leaf_126_wb_clk_i _01899_ _00406_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12492__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15379_ clknet_leaf_125_wb_clk_i _01830_ _00337_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14273__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12952__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold404 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold415 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09940_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] net862 net855 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a22o_1
Xhold459 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09176__A2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09871_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[10\] net722 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__a221o_1
Xfanout917 _04277_ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_2
Xfanout928 net930 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout939 _03421_ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11836__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08822_ net190 net957 _04550_ net1720 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XANTENNA__08923__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10191__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10534__A_N _05257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1126 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net1573 net956 net925 _04533_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
Xhold1148 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07704_ _03593_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nor2_1
XANTENNA__10041__A _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ net747 _04454_ _04466_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07635_ _03492_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14448__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1189_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07566_ _03435_ _03437_ _03456_ team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1
+ vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a211o_1
XANTENNA__09636__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__C _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _04979_ _04980_ _04981_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_1502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09100__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07497_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] team_02_WB.instance_to_wrap.ramload\[8\]
+ net964 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09236_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[25\] net641 net633 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\]
+ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09167_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[27\] net802 net767 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13097__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15531__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14183__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _03993_ _04001_ _03998_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] net823 _04779_ _04780_
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08049_ _03899_ _03935_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold960 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold971 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09167__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold982 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _06247_ _06250_ _06300_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__o31a_1
Xhold993 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[7\] net701 net664 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a22o_1
XANTENNA__11746__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16661__1395 vssd1 vssd1 vccd1 vccd1 net1395 _16661__1395/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16037__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14750_ net1182 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11962_ net344 net2699 net538 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
XANTENNA__09875__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13701_ net1075 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XANTENNA__10485__A1 _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ net911 _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nor2_1
X_14681_ net1193 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XANTENNA__12577__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ net335 net2539 net544 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
X_16420_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[19\]
+ _01294_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13632_ net1071 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10844_ _06401_ _06404_ net366 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16351_ clknet_leaf_96_wb_clk_i _02784_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13563_ net1174 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10775_ net401 _06422_ _06424_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10788__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ clknet_leaf_3_wb_clk_i _01753_ _00260_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12514_ net1805 net321 net479 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16282_ clknet_leaf_101_wb_clk_i _02715_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfxtp_1
XANTENNA__08850__A1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] _03350_ net873 vssd1
+ vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_67_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ clknet_leaf_1_wb_clk_i _01684_ _00191_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12445_ net298 net2264 net484 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XANTENNA__14093__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11510__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09187__A _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ clknet_leaf_63_wb_clk_i _01615_ _00122_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ net273 net1856 net494 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14115_ net1070 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
X_11327_ _06848_ _06941_ net385 vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ clknet_leaf_119_wb_clk_i _01546_ _00053_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09158__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ net1023 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
X_11258_ net434 _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__S net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] net699 net619 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[3\]
+ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08905__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11189_ net410 _06811_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10173__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15997_ clknet_leaf_114_wb_clk_i _02448_ _00955_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14948_ net1034 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XANTENNA__15404__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09330__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14879_ net1162 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
XANTENNA__12487__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16618_ clknet_leaf_61_wb_clk_i _02852_ _01491_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09618__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16549_ clknet_leaf_39_wb_clk_i net1400 _01422_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\] net653 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\]
+ _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09397__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 net132 vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 net140 vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 _02610_ vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 team_02_WB.START_ADDR_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold245 net143 vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 net144 vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 team_02_WB.START_ADDR_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09923_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] net686 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a22o_1
Xfanout703 _04462_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
Xhold289 team_02_WB.instance_to_wrap.top.a1.row1\[104\] vssd1 vssd1 vccd1 vccd1 net1687
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 _04457_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
Xfanout725 _04450_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
XANTENNA_fanout397_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 _04444_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_8
X_09854_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] net872 net832 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a22o_1
Xfanout747 _04440_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10164__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 _04679_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_4
Xfanout769 _04673_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1104_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ net159 net952 net903 net1568 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09785_ _05444_ _05446_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout564_A _07195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08736_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[24\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[24\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08875__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09321__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12397__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\] net702 net698 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout829_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07618_ _03498_ _03504_ _03508_ _03501_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09609__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _04364_ _04373_ _04372_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08607__C team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _03427_ _03438_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ _04764_ _04782_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] net881 net877 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10491_ _05115_ _06034_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ net344 net2170 net514 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ net337 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net521 vssd1
+ vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ net401 _06420_ _06505_ _06738_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12092_ net328 net1980 net526 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold790 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ clknet_leaf_39_wb_clk_i _02371_ _00878_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11043_ _06351_ _06376_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15427__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ clknet_leaf_20_wb_clk_i _02302_ _00809_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_14802_ net1202 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
X_15782_ clknet_leaf_13_wb_clk_i _02233_ _00740_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09848__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11208__C net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _06668_ net226 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ net1035 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11945_ net288 net2271 net536 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14664_ net1008 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
XANTENNA__12100__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net277 net1891 net545 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ clknet_leaf_76_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[2\]
+ _01277_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] sky130_fd_sc_hd__dfrtp_4
X_13615_ net1125 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
X_10827_ _06226_ _06312_ _06474_ net909 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14595_ net1198 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XANTENNA__14816__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16334_ clknet_leaf_100_wb_clk_i _02767_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13546_ net1795 _03383_ net884 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__o21ai_1
X_10758_ net411 _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ clknet_leaf_96_wb_clk_i _00003_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13477_ _03133_ _03309_ _03340_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10689_ team_02_WB.instance_to_wrap.top.pc\[23\] _06340_ vssd1 vssd1 vccd1 vccd1
+ _06341_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15216_ clknet_leaf_34_wb_clk_i _01667_ _00174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ net342 net2365 net489 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__mux2_1
XANTENNA__09379__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16196_ clknet_leaf_66_wb_clk_i _02642_ _01154_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16202__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15147_ clknet_leaf_19_wb_clk_i _01598_ _00105_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12359_ net336 net2187 net496 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15078_ clknet_leaf_59_wb_clk_i _01529_ _00041_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08339__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ net1134 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XANTENNA__10146__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09551__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] net731 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09839__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08521_ net52 net51 net54 net53 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__or4_1
XANTENNA__09303__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12010__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[4\] net917 vssd1 vssd1 vccd1
+ vccd1 _04309_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08383_ _04249_ _04251_ _04252_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16660__1394 vssd1 vssd1 vccd1 vccd1 net1394 _16660__1394/LO sky130_fd_sc_hd__conb_1
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout312_A _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09004_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] net809 net798 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[31\]
+ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09790__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_6
XANTENNA_fanout681_A _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _07216_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_4
Xfanout522 _07212_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09906_ net899 _05548_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o21ai_1
Xfanout533 net535 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09274__B _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_6
Xfanout555 _07198_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_8
Xfanout566 _07195_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_8
X_09837_ _05495_ _05497_ _05499_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__or4_4
Xfanout577 net579 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_4
Xfanout588 _07211_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout946_A _07363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13805__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] net801 net849 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08719_ _04512_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\] net713 net681 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[14\]
+ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08618__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07522__B net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net344 net2454 net564 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11661_ net348 net1723 net573 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
XANTENNA__09058__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _07353_ net995 net940 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__and3b_2
XFILLER_0_119_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10612_ team_02_WB.instance_to_wrap.top.pc\[16\] _06263_ vssd1 vssd1 vccd1 vccd1
+ _06264_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14380_ net1024 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11592_ _06630_ _07177_ _07182_ net438 _07181_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ team_02_WB.instance_to_wrap.top.lcd.nextState\[0\] _03232_ net986 vssd1 vssd1
+ vccd1 vccd1 _03237_ sky130_fd_sc_hd__and3b_1
X_10543_ _05135_ _05153_ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a21oi_2
XANTENNA__16225__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16050_ clknet_leaf_26_wb_clk_i _02501_ _01008_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input75_A wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[4\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[7\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or4_1
X_10474_ _04598_ _04601_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__or2_2
XFILLER_0_126_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15001_ net1190 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12213_ net290 net2567 net512 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12590__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ team_02_WB.START_ADDR_VAL_REG\[1\] net997 net933 vssd1 vssd1 vccd1 vccd1
+ net203 sky130_fd_sc_hd__a21o_1
XANTENNA__09230__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ net274 net2206 net523 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10128__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ net258 net2067 net525 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15903_ clknet_leaf_27_wb_clk_i _02354_ _00861_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11026_ _06144_ _06196_ _06198_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ clknet_leaf_118_wb_clk_i _02285_ _00792_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12977_ _07374_ _07375_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__and2_1
X_15765_ clknet_leaf_115_wb_clk_i _02216_ _00723_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14716_ net1040 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11928_ net346 net2430 net541 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
X_15696_ clknet_leaf_39_wb_clk_i _02147_ _00654_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14647_ net999 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11859_ net333 net2347 net549 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14578_ net1085 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13529_ _03373_ _03374_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16317_ clknet_leaf_80_wb_clk_i _02750_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08272__A2 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16248_ clknet_leaf_92_wb_clk_i _02686_ _01205_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16179_ clknet_leaf_70_wb_clk_i _02625_ _01137_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[14] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_50_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15742__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _03820_ _03823_ net262 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_103_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07883_ _03749_ _03754_ _03756_ _03748_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__or4b_1
XFILLER_0_120_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__S net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[16\] net728 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[16\]
+ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a221o_1
XANTENNA__15892__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[18\] net786 net838 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ team_02_WB.instance_to_wrap.top.a1.hexop\[4\] _04270_ _04326_ vssd1 vssd1
+ vccd1 vccd1 _04336_ sky130_fd_sc_hd__mux2_1
XANTENNA__12292__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] net671 _04499_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XANTENNA__11095__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12796__A_N _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08435_ team_02_WB.instance_to_wrap.top.a1.data\[8\] net916 _04296_ vssd1 vssd1 vccd1
+ vccd1 _04297_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08366_ _04234_ _04235_ _04238_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08799__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08297_ _04154_ _04165_ _04156_ _04155_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15272__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10190_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] net860 net788 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\]
+ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout330 net333 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout341 _03678_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09515__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_4
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
XANTENNA__08723__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
XANTENNA__11754__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ _02927_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__and2b_1
X_13880_ net1055 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XANTENNA__09732__B _05397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ _07375_ _07454_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15550_ clknet_leaf_4_wb_clk_i _02001_ _00508_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12762_ _05175_ _06254_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14501_ net1073 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ net287 net2003 net564 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
X_15481_ clknet_leaf_106_wb_clk_i _01932_ _00439_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12693_ _07257_ _07264_ _07271_ _07291_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12585__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14366__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14432_ net1075 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11644_ net279 net2064 net572 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
X_14363_ net1046 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
Xinput16 wbm_dat_i[18] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ net436 _07166_ _07167_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[1\]
+ sky130_fd_sc_hd__a21o_1
Xinput27 wbm_dat_i[28] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16102_ clknet_leaf_70_wb_clk_i _02548_ _01060_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 wbm_dat_i[9] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ team_02_WB.instance_to_wrap.top.a1.row1\[104\] _03216_ _03219_ team_02_WB.instance_to_wrap.top.a1.row1\[112\]
+ _03213_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__a221o_1
Xinput49 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
XFILLER_0_123_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10526_ _06147_ _06173_ _06175_ _06153_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14294_ net1109 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11929__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16033_ clknet_leaf_2_wb_clk_i _02484_ _00991_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13245_ team_02_WB.instance_to_wrap.ramload\[18\] net980 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[18\] sky130_fd_sc_hd__and2_1
XANTENNA__15765__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13176_ _02781_ _02780_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__nor2_1
X_10388_ _06037_ _06039_ _05032_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__o21a_1
X_12127_ net335 net2001 net586 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09506__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net313 net1871 net530 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11664__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11009_ _05073_ _06037_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15145__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15817_ clknet_leaf_29_wb_clk_i _02268_ _00775_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_16797_ net1351 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
XFILLER_0_90_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15748_ clknet_leaf_55_wb_clk_i _02199_ _00706_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12495__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14276__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ clknet_leaf_27_wb_clk_i _02130_ _00637_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08220_ _04069_ _04101_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08274__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ _04025_ _04032_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08082_ _03950_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11839__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__B _05481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09745__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ _04640_ _04656_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__nor2_4
XFILLER_0_23_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07935_ _03789_ _03794_ _03800_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout477_A _07224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07866_ _03743_ _03755_ _03735_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__a21o_1
XANTENNA__08449__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[17\] net592 vssd1
+ vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__o21ai_2
X_07797_ _03660_ _03671_ net341 _03679_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16070__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout644_A _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13057__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\] net700 net697 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09130__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] net857 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\]
+ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout811_A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08418_ _04268_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__and2b_2
XANTENNA__10291__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09398_ _05052_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15788__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08349_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] _04205_ _04221_ vssd1 vssd1
+ vccd1 vccd1 _04225_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14914__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11360_ _06333_ _06971_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11749__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _05958_ _05960_ _05962_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__or4_2
X_11291_ _06272_ _06278_ _06280_ _04416_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13030_ _07388_ _07389_ _07443_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09197__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] net849 net841 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__a22o_1
XANTENNA__09736__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\] net693 net685 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[4\]
+ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a221o_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1114 net1122 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input38_A wbm_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1205 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_4
Xfanout1158 net1159 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
X_14981_ net1034 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
XANTENNA__13296__A2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1169 net1205 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_2
X_16720_ net1274 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ net1002 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13863_ net1135 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
X_16651_ net1218 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12256__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15602_ clknet_leaf_11_wb_clk_i _02053_ _00560_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12814_ _07396_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16582_ clknet_leaf_82_wb_clk_i net1441 _01455_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13794_ net1088 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12745_ _04764_ _06225_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__or2_1
X_15533_ clknet_leaf_24_wb_clk_i _01984_ _00491_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10282__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15464_ clknet_leaf_56_wb_clk_i _01915_ _00422_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12676_ net420 _06654_ _06901_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14415_ net1112 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11627_ net346 net1734 net577 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
X_15395_ clknet_leaf_45_wb_clk_i _01846_ _00353_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13220__A2 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ net1050 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XANTENNA__10034__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09975__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] net887 net907 team_02_WB.instance_to_wrap.top.pc\[2\]
+ _07151_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11659__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net2006 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ net424 _05836_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__o21ai_1
X_14277_ net1074 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
Xhold619 team_02_WB.instance_to_wrap.top.a1.row2\[2\] vssd1 vssd1 vccd1 vccd1 net2017
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11489_ net426 _07076_ _07079_ _07089_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[5\]
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_29_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16016_ clknet_leaf_39_wb_clk_i _02467_ _00974_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13228_ net1673 net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[1\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09727__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08935__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _03144_ _02784_ _02785_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1308 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1319 team_02_WB.instance_to_wrap.top.a1.row1\[17\] vssd1 vssd1 vccd1 vccd1 net2717
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07720_ _03585_ _03605_ _03609_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13175__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09360__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] _03539_ _03540_ vssd1 vssd1
+ vccd1 vccd1 _03542_ sky130_fd_sc_hd__or3_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07582_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[23\] net686 net634 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15930__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10965__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _04924_ _04926_ _04928_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__or4_4
XFILLER_0_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08203_ _04084_ _04086_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _04857_ _04859_ _04861_ _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13211__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10039__A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08134_ _03981_ _04012_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__xor2_1
XANTENNA__10025__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09966__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08065_ _03932_ _03933_ _03909_ _03925_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1134_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__D _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09179__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09718__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15310__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08878__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _04634_ _04637_ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _03760_ _03808_ _03807_ _03763_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ net459 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09351__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ _03703_ _03737_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14909__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10860_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\] net872 net772 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\]
+ _05176_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a221o_1
X_10791_ _04785_ _06049_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ net1878 net359 net476 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XANTENNA__10264__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_61_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ net343 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[4\] net484 vssd1
+ vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13202__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ net1056 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ _06015_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__and2_1
X_15180_ clknet_leaf_52_wb_clk_i _01631_ _00138_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09957__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12392_ net336 net2116 net494 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08642__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ net1103 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
X_11343_ net301 net2071 net584 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ net1065 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11274_ _05402_ _06024_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13013_ _02958_ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__xnor2_1
X_10225_ _05874_ _05876_ _05878_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__or4_2
XFILLER_0_30_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09590__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\] net871 net791 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[4\]
+ _05799_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[2\] vssd1 vssd1 vccd1 vccd1
+ net1403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12103__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14964_ net1043 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XANTENNA__10412__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09342__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16703_ net1257 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13915_ net1060 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14895_ net1175 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XANTENNA__11942__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16634_ net1382 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
X_13846_ net1084 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07721__A team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16565_ clknet_leaf_99_wb_clk_i net1432 _01438_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13777_ net1028 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
X_10989_ net399 _06622_ _06623_ _06627_ net418 vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15516_ clknet_leaf_62_wb_clk_i _01967_ _00474_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10255__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12728_ _07354_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__inv_2
X_16496_ clknet_leaf_67_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[31\] _01370_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15447_ clknet_leaf_117_wb_clk_i _01898_ _00405_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12659_ _06035_ _06039_ _06044_ _07286_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__A _05296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15378_ clknet_leaf_10_wb_clk_i _01829_ _00336_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ net1063 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
XANTENNA__08081__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold416 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold427 team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] vssd1 vssd1 vccd1 vccd1
+ net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold438 team_02_WB.instance_to_wrap.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net1836
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\] net642 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout907 net908 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
Xfanout918 net920 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout929 net930 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_2
X_08821_ net152 _04341_ _04342_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__o21a_1
XANTENNA__09581__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1116 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[16\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[16\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10322__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1138 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12013__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ _03547_ _03587_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09333__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ net747 _04443_ _04454_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__and3_4
XANTENNA__11852__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _03489_ _03506_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07565_ _03428_ _03432_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout342_A _07116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[24\] net818 net770 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\]
+ _04973_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1084_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07496_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\] team_02_WB.instance_to_wrap.ramload\[9\]
+ net964 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\] net713 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14464__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[27\] net798 net846 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ _03993_ _03998_ _04001_ _03996_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o31a_1
X_09097_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\] net866 net806 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\]
+ _04765_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08048_ _03902_ _03907_ _03932_ _03933_ _03899_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold950 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold972 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold994 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09572__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\] net652 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\]
+ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\] net680 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[7\]
+ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09324__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ net346 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[5\] net538 vssd1
+ vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11762__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ _06343_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__or2_1
X_13700_ net1141 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
X_14680_ net1167 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
XANTENNA__15206__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11892_ net331 net2730 net546 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07541__A team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13631_ net1125 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ _06488_ _06489_ net390 vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11063__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10237__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16350_ clknet_leaf_101_wb_clk_i _02783_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13562_ net1174 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10774_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12513_ net2705 net317 net478 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
X_15301_ clknet_leaf_125_wb_clk_i _01752_ _00259_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16281_ clknet_leaf_94_wb_clk_i _02714_ _01233_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[13\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13493_ _03350_ net873 _03349_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__and3b_1
XANTENNA__12593__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12444_ net288 net1908 net484 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
X_15232_ clknet_leaf_7_wb_clk_i _01683_ _00190_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15163_ clknet_leaf_106_wb_clk_i _01614_ _00121_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12375_ net275 net2721 net493 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__mux2_1
XANTENNA__10945__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14114_ net1093 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11326_ _06895_ _06940_ net380 vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15094_ clknet_leaf_110_wb_clk_i _01545_ _00052_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11937__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ net1105 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
X_11257_ net420 _06124_ _06876_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a21o_1
X_10208_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[3\] net675 net671 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07716__A team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ net418 _06812_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__or2_1
X_10139_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net749 _05796_ vssd1
+ vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__o21a_4
XFILLER_0_94_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15996_ clknet_leaf_48_wb_clk_i _02447_ _00954_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14947_ net1040 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08669__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11672__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ net1191 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16617_ clknet_leaf_60_wb_clk_i _02851_ _01490_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13829_ net1087 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ clknet_leaf_37_wb_clk_i net1438 _01421_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09094__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16479_ clknet_leaf_81_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[14\] _01353_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08841__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09020_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\] net725 net700 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a22o_1
XANTENNA__11701__A team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15849__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08054__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12008__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 team_02_WB.instance_to_wrap.top.a1.data\[10\] vssd1 vssd1 vccd1 vccd1 net1600
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_02_WB.START_ADDR_VAL_REG\[31\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_02_WB.START_ADDR_VAL_REG\[24\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold235 net147 vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 team_02_WB.START_ADDR_VAL_REG\[12\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold257 net120 vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_02_WB.instance_to_wrap.ramload\[28\] vssd1 vssd1 vccd1 vccd1 net1666
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11847__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold279 team_02_WB.instance_to_wrap.top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1 net1677
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[9\] net698 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[9\]
+ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout704 _04461_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 _04457_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09554__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout726 _04450_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_6
X_09853_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] net808 _05506_ _05517_
+ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a211o_1
Xfanout737 _04444_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _04440_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout759 _04679_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout292_A _06935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net160 net951 net902 net1530 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
X_09784_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[12\] net682 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\]
+ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a221o_1
XANTENNA__15229__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ net1591 net958 net924 _04524_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09857__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout557_A _07197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08666_ net748 _04443_ _04446_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08457__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _03503_ _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10872__C1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15379__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ _04383_ _04385_ _04368_ _04378_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout724_A _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16624__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _03435_ _03437_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand2_1
XANTENNA__08607__D team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11967__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07479_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] net2745 net964 vssd1
+ vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08832__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09218_ _04891_ _04893_ _04895_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ _04953_ _06043_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09149_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[27\] net697 net683 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[27\]
+ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__A _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ net334 net2519 net520 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09793__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _05154_ net430 net445 _05155_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__a221o_1
XANTENNA__16004__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15049__RESET_B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ net314 net2153 net526 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold780 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__A1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _05075_ _06663_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__xor2_1
XANTENNA__13257__B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15850_ clknet_leaf_44_wb_clk_i _02301_ _00808_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16154__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A wbm_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14801_ net1199 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
X_15781_ clknet_leaf_128_wb_clk_i _02232_ _00739_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12588__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12993_ _02891_ _02963_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__xnor2_1
X_14732_ net1035 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11944_ net282 net1787 net536 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11875_ net265 net2588 net547 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14663_ net1008 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ clknet_leaf_75_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[1\]
+ _01276_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] sky130_fd_sc_hd__dfrtp_4
X_10826_ _06226_ _06227_ _06311_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__o21bai_1
X_13614_ net1114 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XANTENNA__11407__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__B2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09076__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14594_ net1200 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16333_ clknet_leaf_100_wb_clk_i _02766_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13545_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__and3_1
X_10757_ _06396_ _06407_ net405 vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__mux2_1
XANTENNA__10091__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11521__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13476_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] net2722 vssd1 vssd1 vccd1 vccd1
+ _03340_ sky130_fd_sc_hd__a31o_1
X_16264_ clknet_leaf_101_wb_clk_i _00002_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10688_ team_02_WB.instance_to_wrap.top.pc\[22\] team_02_WB.instance_to_wrap.top.pc\[21\]
+ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15215_ clknet_leaf_33_wb_clk_i _01666_ _00173_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12427_ net348 net2547 net490 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__mux2_1
X_16195_ clknet_leaf_66_wb_clk_i _02641_ _01153_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14832__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09784__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15146_ clknet_leaf_51_wb_clk_i _01597_ _00104_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ net331 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net498 vssd1
+ vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11309_ _05482_ _06021_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__or2_1
X_15077_ clknet_leaf_60_wb_clk_i _01528_ _00040_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12289_ net310 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\] net507 vssd1
+ vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09536__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ net1018 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XANTENNA__09000__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13096__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ clknet_leaf_22_wb_clk_i _02430_ _00937_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ net50 net39 net64 _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08451_ team_02_WB.instance_to_wrap.top.a1.data\[4\] net916 vssd1 vssd1 vccd1 vccd1
+ _04308_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ _04251_ _04252_ _04249_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09067__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15671__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08814__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09003_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] net801 net789 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a22o_1
X_16685__1239 vssd1 vssd1 vccd1 vccd1 _16685__1239/HI net1239 sky130_fd_sc_hd__conb_1
XANTENNA__13034__A1_N _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10909__B1 team_02_WB.instance_to_wrap.top.aluOut\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1047_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15051__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _07218_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09527__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ net897 _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nand2_1
Xfanout512 _07215_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_6
Xfanout523 _07212_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_4
XANTENNA__10137__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_8
XANTENNA_fanout674_A _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net547 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_6
Xfanout556 _07197_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_8
XFILLER_0_67_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09836_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\] net679 net671 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a221o_1
Xfanout567 _07195_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_4
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_6
Xfanout589 _07211_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09767_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\] net821 net785 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[13\]
+ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout841_A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14189__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08718_ _04502_ _04511_ _04514_ _04438_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\] net706 net694 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__and3_2
XFILLER_0_136_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11660_ net339 net2562 net573 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08915__A _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09058__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ net749 _05769_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__o21a_2
XFILLER_0_33_1685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11591_ net423 _06844_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08805__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13330_ team_02_WB.instance_to_wrap.top.a1.row2\[16\] _03234_ _03235_ team_02_WB.instance_to_wrap.top.a1.row2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__a22o_1
X_10542_ _06188_ _06193_ _05156_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ net191 net71 net104 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__and3b_1
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ _04598_ _04601_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nor2_1
XANTENNA__13011__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15000_ net1191 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
X_12212_ net282 net1896 net514 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09766__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ net989 net997 net933 _03173_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__o31a_1
XANTENNA_input68_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__A2 _04908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12143_ net278 net2092 net522 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09518__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ net254 net2316 net525 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
X_15902_ clknet_leaf_3_wb_clk_i _02353_ _00860_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11025_ net450 _06653_ _06661_ net439 _06657_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09481__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__B2 _04527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15833_ clknet_leaf_107_wb_clk_i _02284_ _00791_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11516__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15764_ clknet_leaf_53_wb_clk_i _02215_ _00722_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10420__A _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12111__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15694__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ _02886_ _02965_ net229 vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__o21ai_1
X_14715_ net1033 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ net338 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\] net541 vssd1
+ vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15695_ clknet_leaf_30_wb_clk_i _02146_ _00653_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14827__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10536__A2_N _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14646_ net999 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09049__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11858_ net326 net2392 net549 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10809_ net437 _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11789_ net308 net2674 net559 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14577_ net1080 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ clknet_leaf_96_wb_clk_i _02749_ _01259_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13528_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] _03371_
+ net885 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16247_ clknet_leaf_93_wb_clk_i _02685_ _01204_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_13459_ net1176 _03329_ _03330_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__nor3_1
XANTENNA__15074__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09757__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16178_ clknet_leaf_71_wb_clk_i _02624_ _01136_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_23_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[15] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15129_ clknet_leaf_118_wb_clk_i _01580_ _00087_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 wbm_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09509__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _03821_ _03836_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11316__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07882_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__nor2_2
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__A2 team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[16\] net732 net720 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09552_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[18\] net794 net782 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[18\]
+ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__a221o_1
XANTENNA__12021__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08503_ net2647 _04335_ _04325_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XANTENNA__10827__C1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ _05154_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__and2b_2
XANTENNA__11860__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[8\] net917 vssd1 vssd1 vccd1
+ vccd1 _04296_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08365_ _04227_ _04231_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08799__A1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10055__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08296_ _04168_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout791_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09212__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12704__B _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15567__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08971__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout331 net333 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout342 _07116_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout353 _07153_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
Xfanout364 _05956_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_2
Xfanout375 _05997_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
XANTENNA__09920__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout386 _05909_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
Xfanout397 net398 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_2
X_09819_ _05482_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__and2b_1
X_12830_ _04972_ _06241_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09279__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12740__A_N team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11086__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ _05175_ _06254_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11770__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ net1094 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XANTENNA__10294__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11712_ net279 net1975 net564 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15480_ clknet_leaf_121_wb_clk_i _01931_ _00438_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12692_ _07313_ _07315_ _07319_ _07307_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__o31a_1
X_14431_ net1121 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11643_ net271 net1922 net575 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10046__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09987__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14362_ net1039 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11574_ net449 _07158_ _07165_ net438 _07164_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__a221o_1
Xinput17 wbm_dat_i[19] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 wbm_dat_i[29] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_16101_ clknet_leaf_71_wb_clk_i _02547_ _01059_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput39 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_13313_ _03214_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__nor2_2
X_10525_ _05462_ _05481_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nand2_1
X_14293_ net1121 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ team_02_WB.instance_to_wrap.ramload\[17\] net982 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[17\] sky130_fd_sc_hd__and2_1
XANTENNA__09739__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16032_ clknet_leaf_9_wb_clk_i _02483_ _00990_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ _05883_ net374 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nor2_1
XANTENNA__09203__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13175_ net992 _03150_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__and2_1
XANTENNA__12106__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__A _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _05033_ _06038_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12126_ net332 net2307 net588 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11945__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ net307 net2407 net530 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11701__C_N team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__A2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ net275 net2659 net583 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
XANTENNA__09911__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16684__1238 vssd1 vssd1 vccd1 vccd1 _16684__1238/HI net1238 sky130_fd_sc_hd__conb_1
X_15816_ clknet_leaf_18_wb_clk_i _02267_ _00774_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_16796_ net1350 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
X_15747_ clknet_leaf_40_wb_clk_i _02198_ _00705_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08478__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ _02970_ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11680__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10285__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15678_ clknet_leaf_6_wb_clk_i _02129_ _00636_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14629_ net1157 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10037__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08150_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__inv_2
XANTENNA__09978__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09442__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ team_02_WB.instance_to_wrap.top.a1.row2\[40\] net936 net919 _03968_ vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12805__A _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12016__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08983_ net972 _04632_ _04666_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and3b_4
XANTENNA__11855__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ _03760_ _03820_ _03823_ _03806_ _03809_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a311o_1
X_07865_ _03743_ _03755_ _03735_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _05269_ _05270_ _05272_ _05274_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[17\]
+ sky130_fd_sc_hd__or4_4
X_07796_ _03649_ _03683_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__xor2_2
X_09535_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[18\] net681 net653 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[18\]
+ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout637_A _04488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] net797 net845 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a22o_1
XANTENNA__16365__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08484__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08417_ net919 _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__nor2_1
X_09397_ net897 net612 _04630_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10028__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__inv_2
XANTENNA__10579__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08279_ _04149_ _04150_ _04152_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10310_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[1\] net710 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\]
+ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11290_ _06335_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10241_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[2\] net874 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[2\]
+ _05892_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10200__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10172_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\] net676 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1104 net1138 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
Xfanout1115 net1122 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11765__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1137 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1137 net1138 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
X_14980_ net1041 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_2
X_13931_ net1026 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16650_ net1217 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_13862_ net1142 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15601_ clknet_leaf_16_wb_clk_i _02052_ _00559_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12813_ _05462_ _06276_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__a21o_1
X_16581_ clknet_leaf_67_wb_clk_i net1445 _01454_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13793_ net1102 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10267__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15532_ clknet_leaf_52_wb_clk_i _01983_ _00490_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12744_ _04764_ _06225_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09672__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13205__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ clknet_leaf_16_wb_clk_i _01914_ _00421_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12675_ _06540_ _06634_ net414 vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14414_ net1065 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XANTENNA__11216__C1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11626_ net339 net2583 net577 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
X_15394_ clknet_leaf_47_wb_clk_i _01845_ _00352_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09424__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ net1011 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ team_02_WB.instance_to_wrap.top.pc\[2\] net914 vssd1 vssd1 vccd1 vccd1 _07151_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12625__A _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07719__A team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _05839_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__or2_1
Xhold609 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_2
X_14276_ net1142 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
X_11488_ net434 _07084_ _07085_ net448 _07088_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16015_ clknet_leaf_34_wb_clk_i _02466_ _00973_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ net1686 net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[0\]
+ sky130_fd_sc_hd__and2_1
X_10439_ _06090_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__nand2_1
XANTENNA__14840__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _03148_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__inv_2
XANTENNA__15112__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12109_ net264 net2686 net587 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13089_ team_02_WB.instance_to_wrap.top.pc\[8\] net946 net941 _03099_ vssd1 vssd1
+ vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
Xhold1309 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07650_ _03539_ _03540_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07581_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and2_1
X_16779_ net1333 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_0_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09320_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\] net739 net702 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a22o_1
XANTENNA__10258__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09663__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] net719 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _04011_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__xor2_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[27\] net811 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[27\]
+ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09415__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10039__B team_02_WB.instance_to_wrap.top.DUT.read_data2\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ _03974_ _04002_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07977__A2 _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _03932_ _03933_ _03909_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16799__1353 vssd1 vssd1 vccd1 vccd1 _16799__1353/HI net1353 sky130_fd_sc_hd__conb_1
XFILLER_0_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout587_A _07211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ net886 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15605__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ _03762_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout754_A _04680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net887 _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ _03631_ _03696_ _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__inv_2
XANTENNA__10249__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\] net824 net795 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[19\]
+ _05177_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ net242 net2382 net582 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09654__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[20\] net664 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[20\]
+ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ net347 net2229 net486 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09406__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ _05658_ _05701_ _06014_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12391_ net330 net1964 net494 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14130_ net1082 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
X_11342_ _06887_ _06953_ _06955_ team_02_WB.instance_to_wrap.top.aluOut\[12\] net459
+ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__o32a_2
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16683__1237 vssd1 vssd1 vccd1 vccd1 _16683__1237/HI net1237 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15135__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14061_ net1135 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
X_11273_ _05402_ _06864_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12174__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input50_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] net679 net655 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\]
+ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a221o_1
X_13012_ _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11495__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10155_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] net847 _05811_ _05812_
+ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a211o_1
XANTENNA__15285__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14963_ net1003 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
X_10086_ net899 _05725_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__o21ai_2
Xhold6 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[10\] vssd1 vssd1 vccd1 vccd1
+ net1404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10412__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16702_ net1256 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_13914_ net1058 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14894_ net1175 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ net1381 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
X_13845_ net1120 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16564_ clknet_leaf_82_wb_clk_i net1429 _01437_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13776_ net1021 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
X_10988_ net383 _06483_ net394 vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15515_ clknet_leaf_105_wb_clk_i _01966_ _00473_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12727_ team_02_WB.instance_to_wrap.top.a1.state\[2\] team_02_WB.instance_to_wrap.top.a1.state\[1\]
+ team_02_WB.instance_to_wrap.top.a1.state\[0\] _03419_ vssd1 vssd1 vccd1 vccd1 _07354_
+ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16495_ clknet_leaf_65_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[30\] _01369_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[30\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15446_ clknet_leaf_18_wb_clk_i _01897_ _00404_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ _05236_ _05400_ _06023_ _06029_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11609_ net271 net1995 net579 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__B _05315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15377_ clknet_leaf_18_wb_clk_i _01828_ _00335_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12589_ net333 net2034 net473 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14328_ net1056 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
XANTENNA__08081__A1 team_02_WB.instance_to_wrap.top.a1.row2\[40\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold406 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold417 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16060__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 team_02_WB.instance_to_wrap.top.a1.row1\[15\] vssd1 vssd1 vccd1 vccd1 net1826
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ net1148 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15628__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09030__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12802__B _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout919 net920 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08820_ net153 net954 net903 net1522 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XANTENNA__10191__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1106 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net1580 net957 net925 _04532_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
Xhold1128 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15778__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1139 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10322__B _05975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ _03591_ _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__or2_2
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08682_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\] net670 net667 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a221o_1
XANTENNA__11140__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07633_ _03486_ _03518_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07564_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] _03441_ _03443_ _03451_ vssd1
+ vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__or4_1
XANTENNA__09097__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09636__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09303_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\] net858 net798 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\]
+ _04978_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07495_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] net2749 net964 vssd1
+ vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout335_A _07055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1077_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _04910_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout502_A _07218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08116_ net2592 net936 net919 _04002_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12943__A2 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[29\] net798 net846 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a22o_1
XANTENNA__08072__B2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1352_A team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08047_ _03932_ _03933_ _03908_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_102_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold940 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08889__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold951 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold973 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16553__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold984 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout871_A _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12204__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\] net724 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07583__B1 team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08949_ net972 net886 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13120__A2 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__A_N team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11960_ net339 net2259 net538 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
XANTENNA__09875__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10911_ team_02_WB.instance_to_wrap.top.pc\[26\] _06342_ vssd1 vssd1 vccd1 vccd1
+ _06554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11891_ net326 net2269 net546 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__B team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13630_ net1020 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XANTENNA__09088__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _06394_ _06399_ net366 vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13561_ net1592 net1463 _03395_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08835__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ net580 net401 vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__nand2_2
X_15300_ clknet_leaf_55_wb_clk_i _01751_ _00258_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12512_ net1910 net305 net478 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16280_ clknet_leaf_79_wb_clk_i _02713_ _01232_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13492_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] _03348_ vssd1 vssd1 vccd1
+ vccd1 _03350_ sky130_fd_sc_hd__and2_1
XANTENNA_input98_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ clknet_leaf_27_wb_clk_i _01682_ _00189_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ net281 net2095 net486 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15162_ clknet_leaf_118_wb_clk_i _01613_ _00120_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12374_ net264 net1886 net495 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
XANTENNA__09260__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14113_ net1103 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
X_11325_ _06382_ _06386_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nand2_1
X_15093_ clknet_leaf_115_wb_clk_i _01544_ _00051_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11256_ net580 net420 _06876_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__a21oi_1
X_14044_ net1124 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XANTENNA__09012__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ net897 _05843_ _05861_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o21ai_2
XANTENNA__15920__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _06590_ _06594_ net406 vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__mux2_1
XANTENNA__12114__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ net462 _05769_ _05795_ net456 net740 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a221o_1
X_15995_ clknet_leaf_105_wb_clk_i _02446_ _00953_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11953__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13734__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14946_ net1041 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
X_10069_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\] net787 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[6\]
+ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11122__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09866__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14877_ net1150 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16616_ clknet_leaf_61_wb_clk_i _02850_ _01489_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10881__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ net1142 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09618__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16798__1352 vssd1 vssd1 vccd1 vccd1 _16798__1352/HI net1352 sky130_fd_sc_hd__conb_1
XFILLER_0_134_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16547_ clknet_leaf_0_wb_clk_i net1444 _01420_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ net1118 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XANTENNA__15300__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16478_ clknet_leaf_90_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[13\] _01352_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11701__B _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15429_ clknet_leaf_125_wb_clk_i _01880_ _00387_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15450__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 net121 vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold214 team_02_WB.START_ADDR_VAL_REG\[11\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold225 team_02_WB.instance_to_wrap.top.a1.row1\[121\] vssd1 vssd1 vccd1 vccd1 net1623
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 net134 vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 net133 vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold258 net176 vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 team_02_WB.instance_to_wrap.top.a1.hexop\[2\] vssd1 vssd1 vccd1 vccd1 net1667
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[9\] net702 net673 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09003__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout705 _04461_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
Xfanout716 net719 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_6
XANTENNA__12024__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] net796 net780 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a22o_1
Xfanout727 _04450_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 _04444_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_8
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_2
XANTENNA__10164__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ net161 net953 net905 net1538 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
X_09783_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\] net672 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a22o_1
XANTENNA__11863__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A _06912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08734_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[25\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[25\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10967__A1_N net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ net745 _04445_ _04454_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__and3_1
X_16682__1236 vssd1 vssd1 vccd1 vccd1 _16682__1236/HI net1236 sky130_fd_sc_hd__conb_1
XFILLER_0_7_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1194_A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _03498_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__and2_1
XANTENNA__10872__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _04389_ _04391_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08817__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ _03435_ _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07478_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] net1683 net966 vssd1
+ vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[26\] net863 net807 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[26\]
+ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09148_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\] net706 net677 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _04755_ _04757_ _04759_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__or4_2
XFILLER_0_20_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15943__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12723__A team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ net435 _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net309 net2580 net527 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__mux2_1
Xhold770 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _06037_ _06675_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13341__A2 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10155__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11773__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ net1198 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
X_15780_ clknet_leaf_55_wb_clk_i _02231_ _00738_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12992_ _03012_ _03018_ team_02_WB.instance_to_wrap.top.pc\[24\] net943 vssd1 vssd1
+ vccd1 vccd1 _01522_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09848__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A wbm_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ net1008 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
X_11943_ net274 net1767 net539 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__mux2_1
XANTENNA__11074__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14662_ net1001 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11874_ net259 net1993 net545 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16401_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[0\]
+ _01275_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] sky130_fd_sc_hd__dfrtp_4
X_13613_ net1132 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08808__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10825_ net441 _06440_ _06473_ net428 _06471_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[29\]
+ sky130_fd_sc_hd__a221o_2
X_14593_ net1200 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16332_ clknet_leaf_100_wb_clk_i _02765_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13544_ _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15473__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10756_ _06402_ _06406_ net391 vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16263_ clknet_leaf_96_wb_clk_i _00001_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12109__S net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13475_ _03131_ _03309_ _03339_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10687_ team_02_WB.instance_to_wrap.top.pc\[20\] _06338_ vssd1 vssd1 vccd1 vccd1
+ _06339_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15214_ clknet_leaf_42_wb_clk_i _01665_ _00172_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12426_ net340 net2099 net490 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__mux2_1
X_16194_ clknet_leaf_66_wb_clk_i _02640_ _01152_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11948__S net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ clknet_leaf_29_wb_clk_i _01596_ _00103_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12357_ net327 net2594 net498 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ net449 _06921_ _06924_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__a21oi_1
X_15076_ clknet_leaf_60_wb_clk_i _01527_ _00039_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[29\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ net302 net1984 net505 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08339__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14027_ net1026 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
X_11239_ _06173_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__nand2_1
XANTENNA__10146__A2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11683__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15978_ clknet_leaf_45_wb_clk_i _02429_ _00936_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09839__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14929_ net1000 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08450_ _04307_ net1613 net827 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15816__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08381_ net1760 net935 net918 _04253_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13403__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09472__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12019__S net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\] net767 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09224__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10909__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13639__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ _05567_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[10\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 _07218_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_6
Xfanout513 _07215_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout524 net527 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_6
XFILLER_0_10_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout535 _07206_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_8
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_8
XANTENNA_input5_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] net695 net647 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a22o_1
Xfanout557 _07197_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
Xfanout568 _07193_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_6
Xfanout579 _07189_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout667_A _04478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09766_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\] net814 net841 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13087__B2 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net988 _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout834_A _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] net689 _05364_ vssd1
+ vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15496__CLK clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08579_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12718__A team_02_WB.instance_to_wrap.top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10610_ net929 _05795_ _06220_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09463__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _07178_ _07179_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11270__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ _06188_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13260_ _03174_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.edg2.button_i
+ sky130_fd_sc_hd__inv_2
XANTENNA__09215__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ net420 _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12211_ net274 net1830 net515 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13191_ team_02_WB.START_ADDR_VAL_REG\[0\] _03412_ net932 vssd1 vssd1 vccd1 vccd1
+ _03173_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12142_ net264 net2047 net522 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11069__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16797__1351 vssd1 vssd1 vccd1 vccd1 _16797__1351/HI net1351 sky130_fd_sc_hd__conb_1
X_12073_ net252 net2305 net525 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10128__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11024_ net418 _06658_ _06659_ _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__a22o_1
X_15901_ clknet_leaf_113_wb_clk_i _02352_ _00859_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15832_ clknet_leaf_121_wb_clk_i _02283_ _00790_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15763_ clknet_leaf_3_wb_clk_i _02214_ _00721_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12975_ team_02_WB.instance_to_wrap.top.pc\[26\] net943 net942 _03003_ vssd1 vssd1
+ vccd1 vccd1 _01524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10420__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11008__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14714_ net1042 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
X_11926_ net335 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[7\] net540 vssd1
+ vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
X_15694_ clknet_leaf_40_wb_clk_i _02145_ _00652_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ net999 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11857_ net311 net2515 net549 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
XANTENNA__15989__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11532__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10808_ _06449_ _06456_ net418 vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14576_ net1017 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
X_11788_ net300 net2280 net556 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16315_ clknet_leaf_93_wb_clk_i _02748_ _01258_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_13527_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\] _03371_
+ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__B1 _06880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ _05543_ net370 vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15219__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16246_ clknet_leaf_93_wb_clk_i _02684_ _01203_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[63\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09206__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\]
+ _03326_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11678__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__D team_02_WB.instance_to_wrap.top.aluOut\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12409_ net274 net2715 net490 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__mux2_1
X_16177_ clknet_leaf_71_wb_clk_i _02623_ _01135_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13389_ _03217_ _03221_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__and2b_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11564__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16681__1235 vssd1 vssd1 vccd1 vccd1 _16681__1235/HI net1235 sky130_fd_sc_hd__conb_1
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[26] sky130_fd_sc_hd__buf_2
X_15128_ clknet_leaf_121_wb_clk_i _01579_ _00086_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15369__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07950_ _03831_ _03834_ _03838_ _03839_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a211o_1
X_15059_ clknet_leaf_81_wb_clk_i _01510_ _00022_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10119__A2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07881_ _03767_ _03769_ _03760_ _03762_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09620_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net692 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\]
+ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a221o_1
XANTENNA__12302__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09551_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[18\] net843 net758 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08502_ _02862_ _04326_ _04334_ _04279_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09482_ _05134_ _05153_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09693__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08433_ net960 _04285_ _04294_ _04295_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ _04229_ _04230_ _04227_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__and3b_1
XANTENNA__09445__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08799__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ _04144_ _04159_ _04167_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16144__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11555__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout784_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout310 _06975_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout343 _07116_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout354 net357 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _05956_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net381 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_4
X_09818_ _05461_ _05481_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__nand2_1
Xfanout398 _05863_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12212__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09749_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\] net696 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__a22o_1
XANTENNA__12807__A1 _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ _05134_ _06252_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09684__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11711_ net272 net2050 net566 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ _06796_ _06984_ _07316_ _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__or4_1
XANTENNA__11352__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ net1020 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11642_ net278 net2136 net574 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09436__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ net1059 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
X_11573_ net410 _06819_ _07157_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 wbm_dat_i[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ clknet_leaf_72_wb_clk_i _02546_ _01058_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input80_A wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] team_02_WB.instance_to_wrap.top.lcd.nextState\[4\]
+ _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__or3_2
Xinput29 wbm_dat_i[2] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ _06176_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__inv_2
X_14292_ net1052 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XANTENNA__11498__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16031_ clknet_leaf_26_wb_clk_i _02482_ _00989_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13243_ team_02_WB.instance_to_wrap.ramload\[16\] net982 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[16\] sky130_fd_sc_hd__and2_1
X_10455_ _05929_ net369 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ net992 _03150_ _03151_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _05073_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10415__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output167_A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ net327 net2079 net588 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15661__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ net300 net1754 net530 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11007_ _06641_ _06643_ _06644_ team_02_WB.instance_to_wrap.top.aluOut\[24\] net460
+ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o32a_4
XANTENNA__12122__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15815_ clknet_leaf_16_wb_clk_i _02266_ _00773_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_16795_ net1349 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XANTENNA__16017__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14838__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11961__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15746_ clknet_leaf_51_wb_clk_i _02197_ _00704_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12958_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09675__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ net277 net2037 net542 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ clknet_leaf_117_wb_clk_i _02128_ _00635_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14628_ net1157 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09427__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14559_ net1130 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _03959_ _03965_ _03966_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12982__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15191__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12805__B _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16229_ clknet_leaf_35_wb_clk_i _02674_ _01186_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10606__A team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11537__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ net972 _04632_ _04666_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and3_4
XFILLER_0_80_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07933_ _03760_ _03820_ _03823_ _03809_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_23_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07864_ _03723_ _03732_ _03753_ _03752_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a31o_1
XANTENNA__12032__S net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09603_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] net799 net848 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\]
+ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07795_ team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] _03683_ _03684_ vssd1 vssd1
+ vccd1 vccd1 _03686_ sky130_fd_sc_hd__or3_1
XANTENNA__11871__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _05956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[18\] net725 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09666__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09130__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\] net865 net814 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout532_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08416_ _04271_ _04273_ net916 _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a31o_1
X_16796__1350 vssd1 vssd1 vccd1 vccd1 _16796__1350/HI net1350 sky130_fd_sc_hd__conb_1
X_09396_ net611 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[22\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15534__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ _04208_ _04215_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_102_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _04149_ _04150_ _04152_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout999_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12207__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15684__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[2\] net801 net789 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[2\]
+ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a221o_1
XANTENNA__09197__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[4\] net682 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[4\]
+ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1113 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
Xfanout1116 net1122 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
XFILLER_0_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1127 net1129 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_4
Xfanout1138 net5 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_4
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13930_ net1026 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13861_ net1074 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
X_15600_ clknet_leaf_34_wb_clk_i _02051_ _00558_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11781__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _07400_ _07435_ _07397_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__a21oi_1
X_16580_ clknet_leaf_75_wb_clk_i net1412 _01453_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ net1075 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XANTENNA__09657__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16680__1234 vssd1 vssd1 vccd1 vccd1 _16680__1234/HI net1234 sky130_fd_sc_hd__conb_1
XFILLER_0_70_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15531_ clknet_leaf_19_wb_clk_i _01982_ _00489_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12743_ _04722_ _06222_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15462_ clknet_leaf_11_wb_clk_i _01913_ _00420_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13205__A1 team_02_WB.START_ADDR_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ _06578_ _06605_ net420 vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14413_ net1132 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
X_11625_ _07055_ net2075 net576 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15393_ clknet_leaf_2_wb_clk_i _01844_ _00351_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ net1096 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11556_ _05930_ _06127_ _07150_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[2\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10507_ _06005_ _06159_ _06004_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12117__S net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A3 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14275_ net1069 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XANTENNA__10426__A _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire596 _05790_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_2
X_11487_ net423 net437 _06704_ _07086_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__o311a_1
X_16014_ clknet_leaf_40_wb_clk_i _02465_ _00972_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13226_ _04380_ _04385_ team_02_WB.instance_to_wrap.top.ru.i_ready_i vssd1 vssd1
+ vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.r1.nxt_dmmWen sky130_fd_sc_hd__and3_1
X_10438_ _05461_ net373 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11956__S net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08935__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13157_ _03397_ net895 _03147_ net1183 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a211o_1
X_10369_ _05421_ _05440_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__nor2_1
X_12108_ net261 net1773 net586 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13088_ net890 _07430_ _03096_ _03098_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12039_ net247 net1977 net529 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15407__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09360__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14568__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07580_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] _03438_ vssd1 vssd1 vccd1
+ vccd1 _03471_ sky130_fd_sc_hd__nand2_4
XFILLER_0_125_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08566__A team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778_ net1332 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XFILLER_0_53_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07470__A team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15729_ clknet_leaf_111_wb_clk_i _02180_ _00687_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08320__B1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[25\] net734 net671 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08201_ _04045_ _04047_ _04057_ _04060_ _04046_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__a41o_1
X_09181_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\] net786 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13411__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09820__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08063_ _03940_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__nand2_1
XANTENNA__12027__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09179__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11866__S net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10194__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ net882 _04641_ _04648_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07916_ _03790_ _03791_ _03770_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__a21o_1
X_08896_ _04388_ _04431_ _04433_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__or3_1
XANTENNA__09887__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09860__A _05503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _03696_ _03698_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07778_ _03663_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nor2_1
XANTENNA__09639__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09517_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] net855 _05187_ _05189_
+ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[20\] net704 net676 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13199__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09379_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] net859 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ net426 _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ net328 net1982 net494 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10421__A1 _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11341_ _06276_ net744 _06954_ net913 vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ net1004 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11272_ net267 net2255 net582 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11776__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _07384_ _07386_ _07447_ net888 vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a31o_1
X_10223_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] net711 net635 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[4\] net822 net779 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[4\]
+ _05798_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a221o_1
X_14962_ net1000 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
Xhold7 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[26\] vssd1 vssd1 vccd1 vccd1
+ net1405 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net899 net599 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09342__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ net1255 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_13913_ net1059 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14893_ net1173 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XANTENNA__08550__A0 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13844_ net1052 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
X_16632_ net1380 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_134_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13775_ net1123 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
X_16563_ clknet_leaf_81_wb_clk_i net1450 _01436_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ _06624_ _06625_ net404 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12726_ team_02_WB.instance_to_wrap.top.edg2.flip1 _03403_ _07352_ vssd1 vssd1 vccd1
+ vccd1 _07353_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ clknet_leaf_116_wb_clk_i _01965_ _00472_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16494_ clknet_leaf_65_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[29\] _01368_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ clknet_leaf_115_wb_clk_i _01896_ _00403_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _04742_ _04783_ _04911_ _07284_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ net277 net2298 net578 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ clknet_leaf_37_wb_clk_i _01827_ _00334_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ net326 net2509 net473 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09802__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14327_ net1115 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11539_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[3\] _07119_ vssd1 vssd1 vccd1
+ vccd1 _07135_ sky130_fd_sc_hd__a21o_2
XFILLER_0_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14258_ net1080 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
Xhold429 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11686__S net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13209_ team_02_WB.START_ADDR_VAL_REG\[17\] _04356_ vssd1 vssd1 vccd1 vccd1 net200
+ sky130_fd_sc_hd__and2_1
XFILLER_0_110_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14189_ net1135 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XANTENNA__10176__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout909 _04415_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07465__A team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16355__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08750_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[17\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[17\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__mux2_1
Xhold1107 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07701_ _03548_ net362 _03552_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09333__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08681_ net748 _04442_ _04455_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13406__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _03513_ _03516_ _03520_ _03521_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_36_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12310__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11428__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07563_ team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] _03428_ _03439_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09302_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] net866 net774 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\]
+ _04976_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07494_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] net2742 net965 vssd1
+ vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XANTENNA__10100__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _04888_ _04909_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ _04835_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08115_ _03993_ _03996_ _03998_ _04000_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__o31a_2
X_09095_ _04771_ _04773_ _04775_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08046_ team_02_WB.instance_to_wrap.top.a1.row2\[41\] net936 net920 _03934_ vssd1
+ vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold930 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold952 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold963 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold985 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09572__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09997_ _05656_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout864_A _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15722__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net972 net886 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09324__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08879_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] net916 vssd1 vssd1 vccd1
+ vccd1 _04568_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08918__B _04602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net257 net2578 net585 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XANTENNA__12220__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11890_ net314 net2370 net546 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10841_ _06387_ _06391_ net365 vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13560_ _03360_ _03361_ _03392_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10772_ net413 net396 _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__and3_1
X_12511_ net2301 net297 net476 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15102__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[9\] _03348_ vssd1 vssd1 vccd1
+ vccd1 _03349_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15230_ clknet_leaf_6_wb_clk_i _01681_ _00188_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ net271 net2106 net487 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ clknet_leaf_112_wb_clk_i _01612_ _00119_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12373_ net260 net2395 net495 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15252__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ net1071 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11324_ _06021_ _06938_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__or2_1
X_15092_ clknet_leaf_51_wb_clk_i _01543_ _00050_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14043_ net1061 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11255_ net396 _06650_ _06875_ net409 vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ net897 _05843_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__o21a_1
XANTENNA__09563__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ net407 _06595_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08771__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] _04425_ _05794_ vssd1
+ vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a21o_1
X_15994_ clknet_leaf_123_wb_clk_i _02445_ _00952_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16775__1329 vssd1 vssd1 vccd1 vccd1 _16775__1329/HI net1329 sky130_fd_sc_hd__conb_1
XANTENNA__11658__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14945_ net1043 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\] net815 net791 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12130__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15007__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14876_ net1170 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16615_ clknet_leaf_62_wb_clk_i _02849_ _01488_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_13827_ net1070 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13758_ net1022 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
X_16546_ clknet_leaf_7_wb_clk_i net1454 _01419_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12709_ _05975_ _05936_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__and2b_1
XANTENNA__16483__D team_02_WB.instance_to_wrap.top.aluOut\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13689_ net1064 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16477_ clknet_leaf_81_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[12\] _01351_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15428_ clknet_leaf_18_wb_clk_i _01879_ _00386_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15359_ clknet_leaf_26_wb_clk_i _01810_ _00317_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08054__A2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold204 team_02_WB.START_ADDR_VAL_REG\[22\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold215 team_02_WB.instance_to_wrap.top.a1.row1\[9\] vssd1 vssd1 vccd1 vccd1 net1613
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 team_02_WB.START_ADDR_VAL_REG\[1\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_02_WB.START_ADDR_VAL_REG\[21\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold248 team_02_WB.instance_to_wrap.top.a1.instruction\[0\] vssd1 vssd1 vccd1 vccd1
+ net1646 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[9\] net738 net637 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[9\]
+ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold259 _02609_ vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15745__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12305__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 _04461_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_6
X_09851_ _05510_ _05511_ _05513_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__or4_1
XANTENNA__09554__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 net719 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
Xfanout728 net731 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _04444_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_4
X_08802_ net1625 net953 net904 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09782_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\] net690 _05447_ vssd1
+ vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15895__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ net1608 net958 net924 _04523_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
XANTENNA__09306__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A _06645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12040__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ net746 _04454_ _04455_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__and3_4
X_07615_ _03498_ _03504_ _03505_ _03470_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__a22o_2
XFILLER_0_7_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12799__A_N _05725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10872__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15125__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1187_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _03427_ _03429_ _03433_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net1666 net965 vssd1
+ vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] net851 net787 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16520__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[27\] net674 net653 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\]
+ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09078_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\] net710 net621 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\]
+ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09793__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12723__B team_02_WB.instance_to_wrap.top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08029_ _03914_ _03916_ _03913_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12215__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold760 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold771 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _05075_ _06036_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__nor2_1
Xhold793 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12991_ _04514_ _03015_ _03016_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__and4b_1
XFILLER_0_99_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08648__B team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14730_ net1040 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
X_11942_ net277 net2181 net537 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
XANTENNA__10312__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14661_ net1007 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
X_11873_ net255 net2162 net545 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16400_ clknet_leaf_82_wb_clk_i team_02_WB.instance_to_wrap.top.ru.r1.nxt_dmmRen
+ _01274_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmRen sky130_fd_sc_hd__dfrtp_1
X_13612_ net1004 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
X_10824_ _06212_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nor2_1
XANTENNA__15618__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14592_ net1200 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13543_ net1872 _03381_ net884 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16331_ clknet_leaf_101_wb_clk_i _02764_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10755_ _06404_ _06405_ net366 vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11090__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16262_ clknet_leaf_101_wb_clk_i _00000_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10091__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03339_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10686_ team_02_WB.instance_to_wrap.top.pc\[19\] team_02_WB.instance_to_wrap.top.pc\[18\]
+ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15213_ clknet_leaf_24_wb_clk_i _01664_ _00171_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12425_ net334 net1813 net488 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16193_ clknet_leaf_65_wb_clk_i _02639_ _01151_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15144_ clknet_leaf_55_wb_clk_i _01595_ _00102_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12356_ net311 net2287 net498 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__mux2_1
XANTENNA__09784__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _06022_ net432 _06922_ net438 _06923_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__a221o_1
X_15075_ clknet_leaf_60_wb_clk_i _01526_ _00038_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[28\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12125__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__A _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ net293 net2465 net504 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14026_ net1050 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XANTENNA__09536__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _06174_ _06858_ _05572_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__a21o_1
XANTENNA__11964__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ net417 _06795_ _06412_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15148__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15977_ clknet_leaf_24_wb_clk_i _02428_ _00935_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14928_ net1001 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10303__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14859_ net1174 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15298__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _04251_ _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold99_A team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16529_ clknet_leaf_75_wb_clk_i team_02_WB.instance_to_wrap.top.ru.i_ready_i _01403_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.i_ready sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07483__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10082__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[31\] net813 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12035__S net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09527__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09903_ _05557_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 _07218_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout514 _07215_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_8
Xfanout525 net527 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08735__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11334__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 net539 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_8
Xfanout547 _07201_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_4
X_09834_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\] net707 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[11\]
+ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1102_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _07193_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_4
X_09765_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\] net765 _05431_ vssd1
+ vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16073__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11175__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__B _04277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _04360_ net463 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__or2_1
X_09696_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] net662 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a22o_1
XANTENNA__09160__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ net746 _04442_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and3_4
XFILLER_0_7_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ _04370_ net978 net979 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or3b_2
XFILLER_0_33_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07529_ team_02_WB.instance_to_wrap.top.a1.state\[2\] _03420_ vssd1 vssd1 vccd1 vccd1
+ _03422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15910__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07474__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ _06184_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__or2_1
XANTENNA__11270__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16774__1328 vssd1 vssd1 vccd1 vccd1 _16774__1328/HI net1328 sky130_fd_sc_hd__conb_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ net396 _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12210_ net275 net2493 net513 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13190_ _02785_ _03162_ _03171_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o21a_1
XANTENNA__09766__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12141_ net260 net2035 net523 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09518__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ net247 net1855 net525 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold590 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11784__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ clknet_leaf_63_wb_clk_i _02351_ _00858_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16416__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net394 _06072_ net416 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13565__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15831_ clknet_leaf_119_wb_clk_i _02282_ _00789_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12974_ _06555_ _07336_ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__o21ai_1
X_15762_ clknet_leaf_25_wb_clk_i _02213_ _00720_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1290 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
X_14713_ net1042 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11925_ net330 net2183 net541 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XANTENNA_output112_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15693_ clknet_leaf_32_wb_clk_i _02144_ _00651_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ net307 net2087 net551 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
X_14644_ net1002 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12628__B _06846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _06452_ _06455_ net407 vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__mux2_1
X_14575_ net1129 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10429__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15590__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ net293 net2714 net556 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
X_16314_ clknet_leaf_77_wb_clk_i _02747_ _01257_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13526_ _03371_ _03372_ net885 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__and3b_1
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10738_ _05591_ net375 vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__S net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13457_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] _03326_ net1653 vssd1
+ vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16245_ clknet_leaf_93_wb_clk_i _02683_ _01202_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ net581 _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ net275 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[24\] net489 vssd1
+ vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09757__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16176_ clknet_leaf_71_wb_clk_i _02622_ _01134_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_13388_ net2405 net896 _03288_ net993 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__o211a_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_2_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[17] sky130_fd_sc_hd__buf_2
X_12339_ net256 net2485 net499 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
X_15127_ clknet_leaf_117_wb_clk_i _01578_ _00085_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_107_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08983__A_N net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09509__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15058_ clknet_leaf_91_wb_clk_i _01509_ _00021_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11694__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ net1062 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07880_ _03763_ _03770_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08569__A team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09550_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[18\] net806 net767 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\]
+ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08501_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] net990 _04276_ vssd1 vssd1
+ vccd1 vccd1 _04334_ sky130_fd_sc_hd__or3_1
X_09481_ _05134_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15933__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ net2717 net827 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ _04235_ _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10055__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08294_ _04106_ _04132_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11869__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout310_A _06975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout408_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12201__B1 _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07759__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15313__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08971__A3 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 net302 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
Xfanout311 _06996_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11307__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 _06834_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
Xfanout333 _07035_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout344 _07116_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
Xfanout355 net357 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12720__C team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 _05956_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_2
XANTENNA__09381__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 net381 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09920__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _05461_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__nor2_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_2
XANTENNA_fanout944_A _07363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout399 net402 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09748_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\] net688 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\]
+ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[15\] net857 net789 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[15\]
+ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a221o_1
XANTENNA__11633__A team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ net275 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[24\] net566 vssd1
+ vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10294__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ _06684_ _06823_ _06851_ _07317_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11641_ net264 net2638 net575 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14360_ net1105 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XANTENNA__10046__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ net422 _06811_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__nor2_1
XANTENNA__09987__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13311_ net986 net987 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__or2_2
XANTENNA__11779__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 wbm_dat_i[20] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ _05421_ _05440_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__and2b_1
X_14291_ net1149 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
X_13242_ net1647 net983 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmload_co\[15\]
+ sky130_fd_sc_hd__and2_1
X_16030_ clknet_leaf_3_wb_clk_i _02481_ _00988_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10454_ _06104_ _06106_ net365 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input73_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13173_ _03148_ _03159_ _03160_ _03149_ _03157_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a32o_1
X_10385_ _05012_ _05030_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12124_ net313 net2507 net588 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__mux2_1
XANTENNA__15806__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12055_ net292 net1939 net528 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XANTENNA__12403__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _06242_ net743 net457 team_02_WB.instance_to_wrap.top.a1.dataIn\[24\] net443
+ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__a221o_1
XANTENNA__09372__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15814_ clknet_leaf_3_wb_clk_i _02265_ _00772_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_16794_ net1348 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XANTENNA__09124__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15745_ clknet_leaf_3_wb_clk_i _02196_ _00703_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12957_ _07366_ _02985_ _02988_ _07364_ team_02_WB.instance_to_wrap.top.pc\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__o32a_1
XFILLER_0_38_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08478__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11908_ net264 net1968 net542 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10285__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15676_ clknet_leaf_61_wb_clk_i _02127_ _00634_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12888_ team_02_WB.instance_to_wrap.top.pc\[6\] _05771_ vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14627_ net1156 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
X_11839_ net252 net2090 net550 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10037__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11234__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09978__A2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14558_ net1020 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11689__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12982__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _03359_ _03360_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\] vssd1 vssd1 vccd1
+ vccd1 _03361_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16491__D team_02_WB.instance_to_wrap.top.aluOut\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14489_ net1064 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16228_ clknet_leaf_35_wb_clk_i _02673_ _01185_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07468__A team_02_WB.instance_to_wrap.top.a1.dataIn\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12734__A1 _07352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07940__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16159_ clknet_leaf_35_wb_clk_i net1495 _01117_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15486__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _04637_ _04641_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07932_ _03821_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__and2_1
XANTENNA__13409__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07863_ _03723_ _03732_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09602_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[17\] net867 net881 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a22o_1
X_16773__1327 vssd1 vssd1 vccd1 vccd1 _16773__1327/HI net1327 sky130_fd_sc_hd__conb_1
X_07794_ _03683_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__or2_1
XANTENNA__09115__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ _05198_ _05200_ _05202_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__or4_4
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\] net801 net849 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\]
+ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a221o_1
XANTENNA__11473__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ _04279_ _04280_ _04281_ net937 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a22o_1
X_09395_ _05064_ _05068_ _05069_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__nor4_2
XANTENNA_fanout525_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10028__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A _05503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _04204_ _04218_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nor2_1
XANTENNA__09969__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08277_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04153_ _04155_ _04156_ vssd1
+ vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_127_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15829__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10200__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10170_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[4\] net672 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1106 net1113 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
Xfanout1117 net1122 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12223__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_2
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15209__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860_ net1142 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09106__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ _07399_ _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ net1130 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ clknet_leaf_44_wb_clk_i _01981_ _00488_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10267__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12742_ net988 team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1 _07366_
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_112_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15461_ clknet_leaf_128_wb_clk_i _01912_ _00419_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12673_ net414 _06506_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13205__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16604__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__A2 _04315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11216__A1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14412_ net1012 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
X_11624_ net333 net1906 net577 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15392_ clknet_leaf_10_wb_clk_i _01843_ _00350_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12906__B _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ net1136 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
X_11555_ net448 _07141_ _07146_ net434 _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10707__A _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10506_ net386 _05929_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14274_ net1091 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_11486_ _06011_ net454 vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12716__A1 team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10426__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire597 _05790_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_2
X_13225_ _04374_ team_02_WB.instance_to_wrap.top.ru.i_ready_i vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.r1.nxt_dmmRen sky130_fd_sc_hd__and2_1
X_16013_ clknet_leaf_21_wb_clk_i _02464_ _00971_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10437_ _05421_ net367 vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09593__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13156_ team_02_WB.instance_to_wrap.top.lcd.currentState\[5\] net895 vssd1 vssd1
+ vccd1 vccd1 _03147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ _05484_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ net256 net2595 net589 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10442__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _07032_ net227 _03097_ net230 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12133__S net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ _05939_ _05947_ _05951_ _05953_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[1\]
+ sky130_fd_sc_hd__or4_4
XANTENNA__09345__B1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ net245 net1824 net529 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11972__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16134__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16486__D team_02_WB.instance_to_wrap.top.aluOut\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16777_ net1331 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
X_13989_ net1087 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XANTENNA__08566__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15728_ clknet_leaf_42_wb_clk_i _02179_ _00686_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10258__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15659_ clknet_leaf_21_wb_clk_i _02110_ _00617_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08200_ _04041_ _04061_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12404__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\] net771 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08131_ _03944_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12308__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ _03945_ _03946_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09584__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A team_02_WB.instance_to_wrap.top.a1.dataIn\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12043__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] _04643_ vssd1 vssd1
+ vccd1 vccd1 _04649_ sky130_fd_sc_hd__or2_1
XANTENNA__10352__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1015_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09336__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ _03779_ _03804_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__or3b_1
X_08895_ net594 _04578_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11882__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07846_ _03710_ _03715_ _03717_ _03708_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09860__B _05521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07777_ _03621_ _03645_ _03632_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15501__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\] net804 net784 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[19\]
+ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a221o_1
XANTENNA__10249__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11446__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09447_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] net701 _05120_ vssd1
+ vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09378_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\] net814 net775 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a22o_1
XANTENNA__15651__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08329_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04165_ vssd1 vssd1 vccd1
+ vccd1 _04206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12218__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ team_02_WB.instance_to_wrap.top.pc\[12\] _06333_ vssd1 vssd1 vccd1 vccd1
+ _06954_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10421__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13032__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16007__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ _06885_ _06887_ _06890_ team_02_WB.instance_to_wrap.top.aluOut\[15\] net461
+ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__o32a_4
XANTENNA__12742__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ team_02_WB.instance_to_wrap.top.pc\[21\] net944 net941 _03033_ vssd1 vssd1
+ vccd1 vccd1 _01519_ sky130_fd_sc_hd__a22o_1
XANTENNA__09575__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\] net731 net723 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\]
+ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a221o_1
XANTENNA__07836__A team_02_WB.instance_to_wrap.top.a1.dataIn\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\] net811 net851 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16157__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A wbm_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net598 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[6\]
+ sky130_fd_sc_hd__inv_2
X_14961_ net1001 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XANTENNA__11792__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[21\] vssd1 vssd1 vccd1 vccd1
+ net1406 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ net1254 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13573__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ net1057 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14892_ net1173 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16631_ net1379 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15181__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ net1148 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16562_ clknet_leaf_39_wb_clk_i net1460 _01435_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13774_ net1116 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
X_10986_ net386 _06492_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15513_ clknet_leaf_106_wb_clk_i _01964_ _00471_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12725_ _04359_ _07346_ _07349_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__and4b_2
X_16493_ clknet_leaf_65_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[28\] _01367_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08853__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15444_ clknet_leaf_53_wb_clk_i _01895_ _00402_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _04699_ _04824_ _05524_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ net263 net2237 net578 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15375_ clknet_leaf_35_wb_clk_i _01826_ _00333_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12128__S net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12587_ net311 net2667 net473 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA__10437__A _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14326_ net1110 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16772__1326 vssd1 vssd1 vccd1 vccd1 _16772__1326/HI net1326 sky130_fd_sc_hd__conb_1
X_11538_ _07131_ _07132_ _07134_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[3\]
+ sky130_fd_sc_hd__or3_2
XFILLER_0_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold408 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold419 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _05747_ net432 _07057_ _07071_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[6\]
+ sky130_fd_sc_hd__a211o_1
X_14257_ net1029 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13208_ team_02_WB.START_ADDR_VAL_REG\[16\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net199 sky130_fd_sc_hd__a21o_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09030__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188_ net1004 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
X_13139_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[3\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__and4_1
XANTENNA__09318__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15524__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14579__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _03548_ _03552_ net362 vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08680_ net745 _04446_ _04455_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__and3_4
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07631_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07562_ _03441_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15674__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\] net875 net754 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\]
+ _04977_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07493_ team_02_WB.instance_to_wrap.top.a1.instruction\[12\] team_02_WB.instance_to_wrap.ramload\[12\]
+ net969 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08844__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ _04869_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ _04837_ _04839_ _04841_ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__or4_1
XANTENNA__12038__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13050__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08114_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09094_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] net790 net838 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[29\]
+ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11877__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ _03932_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold920 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold931 team_02_WB.instance_to_wrap.top.pad.keyCode\[4\] vssd1 vssd1 vccd1 vccd1
+ net2329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09557__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13353__B2 team_02_WB.instance_to_wrap.top.a1.row2\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold953 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09021__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold964 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold975 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold986 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09996_ _05633_ _05655_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__and2_1
XANTENNA__09309__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net977 _04369_ _04368_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12501__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08878_ net1556 _04567_ net825 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
X_07829_ _03682_ _03686_ _03687_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10840_ net363 _06350_ _06351_ _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__a31o_1
XANTENNA__11419__A1 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09088__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ _06417_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08835__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16719__1273 vssd1 vssd1 vccd1 vccd1 _16719__1273/HI net1273 sky130_fd_sc_hd__conb_1
XFILLER_0_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12510_ net2221 net289 net476 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ _03348_ net873 _03347_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__and3b_1
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net276 net2510 net485 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14952__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12372_ net254 net1835 net493 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__mux2_1
X_15160_ clknet_leaf_122_wb_clk_i _01611_ _00118_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09260__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__A team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14111_ net1130 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
X_11323_ _05484_ _06020_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__nor2_1
XANTENNA__11787__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15091_ clknet_leaf_126_wb_clk_i _01542_ _00049_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09548__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14042_ net1052 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
X_11254_ net393 _06874_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__nand2_1
XANTENNA__09012__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[3\] vssd1 vssd1 vccd1
+ vccd1 _05861_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11185_ net427 _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16629__1377 vssd1 vssd1 vccd1 vccd1 net1377 _16629__1377/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08771__B2 _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04367_ _04426_ net972
+ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15993_ clknet_leaf_117_wb_clk_i _02444_ _00951_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10067_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[6\] net880 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a22o_1
XANTENNA__12411__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14944_ net1008 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XANTENNA__10720__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875_ net1190 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16614_ clknet_leaf_57_wb_clk_i _02848_ _01487_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ net1088 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16545_ clknet_leaf_28_wb_clk_i net1416 _01418_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13757_ net1031 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10969_ net441 _06588_ _06589_ net428 vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10094__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ _04513_ _07335_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16476_ clknet_leaf_91_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[11\] _01350_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[11\] sky130_fd_sc_hd__dfrtp_1
X_13688_ net1107 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15427_ clknet_leaf_45_wb_clk_i _01878_ _00385_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13032__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ _04744_ _04785_ _07266_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14862__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15077__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09787__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15358_ clknet_leaf_4_wb_clk_i _01809_ _00316_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09251__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11697__S net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold205 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] vssd1
+ vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ net1073 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
Xhold216 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] vssd1 vssd1
+ vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ clknet_leaf_112_wb_clk_i _01740_ _00247_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold227 net162 vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 team_02_WB.START_ADDR_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 team_02_WB.instance_to_wrap.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net1647
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09003__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16472__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[11\] net803 net768 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[11\]
+ _05514_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout707 _04461_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 net731 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ net163 net953 net904 net1512 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a22o_1
X_09781_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\] net704 net698 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a22o_1
XANTENNA__13099__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08732_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[26\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[26\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XANTENNA__12321__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08663_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] net723 net719 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\]
+ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ team_02_WB.instance_to_wrap.top.a1.dataIn\[30\] _03438_ _03499_ vssd1 vssd1
+ vccd1 vccd1 _03505_ sky130_fd_sc_hd__a21o_1
XANTENNA__10872__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08594_ net976 _04377_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ _03431_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1
+ _03436_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08817__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_A _07075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1082_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07476_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] net1707 net965 vssd1
+ vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09490__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\] net800 net762 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\]
+ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[27\] net717 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09778__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[29\] net669 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__inv_2
XANTENNA__12723__C team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold750 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold761 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold783 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08753__B2 _04533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09979_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] net795 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[8\]
+ _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a221o_1
XANTENNA__10560__A1 _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12990_ _07376_ _07377_ _07452_ _07453_ net888 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a311o_1
XFILLER_0_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09702__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11941_ net263 net2603 net537 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16771__1325 vssd1 vssd1 vccd1 vccd1 _16771__1325/HI net1325 sky130_fd_sc_hd__conb_1
XFILLER_0_19_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14660_ net1000 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11872_ net253 net2085 net545 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_1
XANTENNA__08945__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13611_ net1026 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
X_10823_ _04785_ _06211_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08808__A2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14591_ net1200 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ clknet_leaf_100_wb_clk_i _02763_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13542_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\] _03381_
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16345__CLK clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ _04502_ net374 vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16261_ clknet_leaf_93_wb_clk_i _02699_ _01218_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[109\]
+ sky130_fd_sc_hd__dfstp_1
X_10685_ team_02_WB.instance_to_wrap.top.pc\[17\] _06336_ vssd1 vssd1 vccd1 vccd1
+ _06337_ sky130_fd_sc_hd__and2_1
X_13473_ _03130_ _03309_ _03338_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15212_ clknet_leaf_52_wb_clk_i _01663_ _00170_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09769__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ net331 net2738 net490 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__mux2_1
X_16192_ clknet_leaf_64_wb_clk_i _02638_ _01150_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ clknet_leaf_15_wb_clk_i _01594_ _00101_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_12355_ net309 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[11\] net498 vssd1
+ vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__mux2_1
XANTENNA__12406__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10715__A _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11306_ _05441_ net446 _06149_ net454 vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__a22o_1
X_15074_ clknet_leaf_60_wb_clk_i _01525_ _00037_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12286_ net286 net1742 net506 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__mux2_1
XANTENNA__10434__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14025_ net1024 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
X_11237_ _06146_ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10000__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09941__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ net407 _06566_ _06567_ _06793_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[5\] net819 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[5\]
+ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12141__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10450__A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ _05156_ _06194_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15976_ clknet_leaf_85_wb_clk_i _02427_ _00934_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09016__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14927_ net999 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11980__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13761__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14858_ net1174 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16494__D team_02_WB.instance_to_wrap.top.aluOut\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ net1028 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14789_ net1177 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10067__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ clknet_leaf_39_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[31\]
+ _01402_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09472__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16459_ clknet_leaf_58_wb_clk_i net1542 _01333_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09000_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\] net782 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ _04684_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09224__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12316__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13001__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09902_ _05559_ _05561_ _05563_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12840__A _04624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 net507 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_6
Xfanout515 _07215_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16718__1272 vssd1 vssd1 vccd1 vccd1 _16718__1272/HI net1272 sky130_fd_sc_hd__conb_1
XANTENNA__08735__B2 _04524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_8
X_09833_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[11\] net735 net691 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a22o_1
Xfanout537 net539 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_8
Xfanout548 _07200_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_6
Xfanout559 _07197_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_4
XANTENNA__10542__A1 _06188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A _06727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09764_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\] net878 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08715_ _04502_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__nor2_1
X_09695_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\] net677 net669 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\]
+ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11890__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_136_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15242__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__and3_2
XFILLER_0_90_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16638__1209 vssd1 vssd1 vccd1 vccd1 _16638__1209/HI net1209 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08577_ _04364_ _04371_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout722_A _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10058__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12718__C team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09999__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ team_02_WB.instance_to_wrap.top.a1.state\[2\] _03420_ vssd1 vssd1 vccd1 vccd1
+ _03421_ sky130_fd_sc_hd__and2_1
XANTENNA__09463__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16628__1376 vssd1 vssd1 vccd1 vccd1 net1376 _16628__1376/LO sky130_fd_sc_hd__conb_1
XFILLER_0_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ team_02_WB.instance_to_wrap.top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 _03400_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11270__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ net388 _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09215__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09129_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[28\] net794 net875 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[28\]
+ _04806_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a221o_1
XANTENNA__12226__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ net257 net2102 net522 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10781__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net244 net2207 net525 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12750__A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold580 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ net399 _06101_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__nand2_1
XANTENNA__09923__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15830_ clknet_leaf_110_wb_clk_i _02281_ _00788_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15761_ clknet_leaf_16_wb_clk_i _02212_ _00719_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12973_ net229 _03000_ _03001_ _02866_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_38_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1280 team_02_WB.instance_to_wrap.ramload\[8\] vssd1 vssd1 vccd1 vccd1 net2678
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ net1008 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10297__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13581__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ net327 net2709 net541 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
X_15692_ clknet_leaf_52_wb_clk_i _02143_ _00650_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14643_ net1040 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11855_ net299 net2138 net548 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10806_ _06453_ _06454_ net391 vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__mux2_1
X_14574_ net1116 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
X_11786_ net285 net1987 net558 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XANTENNA__09454__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10429__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16313_ clknet_leaf_80_wb_clk_i _02746_ _01256_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13525_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\]
+ _03366_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] vssd1
+ vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10737_ _06384_ _06387_ net365 vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__mux2_1
XANTENNA__11261__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16244_ clknet_leaf_93_wb_clk_i _02682_ _01201_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13456_ net2006 _03326_ _03328_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10668_ _04431_ _04433_ _04388_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__or3b_1
XANTENNA__09206__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ net263 net2077 net489 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16175_ clknet_leaf_66_wb_clk_i _02621_ _01133_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12136__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__A _05633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ _03287_ _03206_ _03277_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__or3b_1
X_10599_ team_02_WB.instance_to_wrap.top.pc\[21\] _06248_ vssd1 vssd1 vccd1 vccd1
+ _06251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10221__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
X_15126_ clknet_leaf_111_wb_clk_i _01577_ _00084_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 wbm_adr_o[18] sky130_fd_sc_hd__buf_2
X_12338_ net253 net1938 net497 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11975__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15057_ clknet_leaf_91_wb_clk_i _01508_ _00020_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_12269_ net239 net2737 net506 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14008_ net1057 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XANTENNA__09914__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16489__D team_02_WB.instance_to_wrap.top.aluOut\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07473__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16510__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ clknet_leaf_119_wb_clk_i _02410_ _00917_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09142__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ net1798 _04332_ _04325_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XANTENNA__10288__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09480_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[20\] net592 vssd1
+ vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09693__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ team_02_WB.instance_to_wrap.top.a1.data\[9\] net915 _04293_ vssd1 vssd1 vccd1
+ vccd1 _04294_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08362_ net1685 net935 net918 _04236_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08658__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09445__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08293_ _04170_ _04171_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12046__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _06780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16770__1324 vssd1 vssd1 vccd1 vccd1 _16770__1324/HI net1324 sky130_fd_sc_hd__conb_1
XANTENNA__10212__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11885__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16040__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
Xfanout312 _06996_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15608__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 net325 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout672_A _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _07116_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_1
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12720__D team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_2
X_09816_ net897 _05480_ _04630_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a21o_1
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_2
Xfanout389 _05908_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16190__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09747_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[13\] net712 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15758__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[15\] net793 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a22o_1
XANTENNA__09684__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__B _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ net977 _04370_ net889 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11640_ net258 net2020 net572 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09436__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ net429 _06156_ _07161_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12745__A _04764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13310_ _03214_ _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__nor2_2
XFILLER_0_68_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ _05633_ _05655_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__nand2b_1
X_14290_ net1081 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15138__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13241_ team_02_WB.instance_to_wrap.ramload\[14\] net983 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[14\] sky130_fd_sc_hd__and2_1
X_10453_ _05836_ net374 _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10203__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input66_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13172_ _03154_ _03156_ _03158_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o21ai_1
X_10384_ _05075_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11795__S net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ net309 net2228 net589 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13576__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15288__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12054_ net283 net2429 net529 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XANTENNA__10506__A1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11005_ net911 _06642_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nor2_1
X_15813_ clknet_leaf_127_wb_clk_i _02264_ _00771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout890 _04362_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_4
X_16793_ net1347 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_0_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15744_ clknet_leaf_11_wb_clk_i _02195_ _00702_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12956_ _02972_ _02984_ _02987_ _04362_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07513__S _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11907_ net258 net1942 net542 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15675_ clknet_leaf_106_wb_clk_i _02126_ _00633_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12887_ team_02_WB.instance_to_wrap.top.pc\[6\] _05771_ vssd1 vssd1 vccd1 vccd1 _02921_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14626_ net1156 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11838_ net247 net2426 net550 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09427__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16717__1271 vssd1 vssd1 vccd1 vccd1 _16717__1271/HI net1271 sky130_fd_sc_hd__conb_1
XFILLER_0_83_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11234__A2 team_02_WB.instance_to_wrap.top.aluOut\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14557_ net1054 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
X_11769_ net240 net2623 net558 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15031__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__or4_1
XANTENNA__07989__A2 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12982__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14488_ net1062 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16227_ clknet_leaf_30_wb_clk_i _02672_ _01184_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13439_ _03303_ _03307_ net1678 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16158_ clknet_leaf_37_wb_clk_i net1511 _01116_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16637__1208 vssd1 vssd1 vccd1 vccd1 _16637__1208/HI net1208 sky130_fd_sc_hd__conb_1
XFILLER_0_122_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15109_ clknet_leaf_128_wb_clk_i _01560_ _00067_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _04634_ _04636_ _04637_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and3_1
X_16089_ clknet_leaf_80_wb_clk_i _02535_ _01047_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ _03769_ _03810_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15900__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _03713_ _03745_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__xnor2_4
X_09601_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[17\] net872 net815 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\]
+ _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a221o_1
X_07793_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] net341 _03679_ vssd1 vssd1
+ vccd1 vccd1 _03684_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[18\] net729 net669 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[18\]
+ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a221o_1
XANTENNA__09666__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09463_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\] net761 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout253_A _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ _04268_ net961 vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__nor2_1
X_09394_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] net819 net811 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\]
+ _05055_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08345_ _04207_ _04215_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__xor2_1
XANTENNA__12565__A team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B _05521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13160__S _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ _04146_ _04152_ _04148_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10085__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16556__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12504__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1107 net1113 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_4
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
Xfanout1129 net1137 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15580__CLK clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _05544_ _05548_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14020__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13790_ net1022 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09657__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net988 team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1 _07365_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_96_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15460_ clknet_leaf_54_wb_clk_i _01911_ _00418_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12672_ net414 _06418_ _06468_ net435 _06125_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14411_ net1027 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
X_11623_ net329 net2066 net577 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
X_15391_ clknet_leaf_26_wb_clk_i _01842_ _00349_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ net1147 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
X_11554_ net423 net437 _06797_ _07148_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__o31a_1
XFILLER_0_110_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09290__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ _05934_ _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__and2b_1
X_14273_ net1145 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11485_ _05793_ net432 _06135_ _06009_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_46_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16012_ clknet_leaf_23_wb_clk_i _02463_ _00970_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13224_ team_02_WB.instance_to_wrap.busy_o net968 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.i_ready_i
+ sky130_fd_sc_hd__and2b_1
Xwire598 net600 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09042__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08396__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15923__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ _03146_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__inv_2
XANTENNA__12414__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__A _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ _05522_ _06019_ _05524_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a21o_1
X_12106_ net251 net2415 net587 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13086_ _02917_ _02938_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__xor2_1
X_10298_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[1\] net817 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[1\]
+ _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12037_ net237 net1928 net529 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11152__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16776_ net1330 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13988_ net1141 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
X_15727_ clknet_leaf_31_wb_clk_i _02178_ _00685_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08856__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ team_02_WB.instance_to_wrap.top.pc\[29\] _06229_ _02972_ vssd1 vssd1 vccd1
+ vccd1 _02973_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16429__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08320__A2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15658_ clknet_leaf_44_wb_clk_i _02109_ _00616_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14609_ net1196 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15589_ clknet_leaf_128_wb_clk_i _02040_ _00547_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] _03967_ vssd1 vssd1 vccd1
+ vccd1 _04016_ sky130_fd_sc_hd__or2_2
XFILLER_0_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09820__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ _03906_ _03934_ _03938_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12324__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] _04643_ vssd1 vssd1
+ vccd1 vccd1 _04648_ sky130_fd_sc_hd__nor2_2
XANTENNA__10352__B _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ _03780_ _03795_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nand2_2
XANTENNA__12340__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09887__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07845_ _03710_ _03715_ _03717_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout370_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout468_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07776_ _03617_ _03655_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__xor2_2
XANTENNA__09639__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\] net864 net808 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08847__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09446_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[20\] net624 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13199__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout802_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ _05052_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ _04202_ _04203_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09811__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15946__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _04127_ _04130_ _04134_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09024__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ _06266_ net743 _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _06889_
+ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a221o_1
XANTENNA__12742__B team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] net719 net703 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12234__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10152_ _05803_ _05805_ _05807_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__or4_1
X_14960_ net999 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
X_10083_ _05736_ _05740_ _05741_ _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__nor4_2
X_16716__1270 vssd1 vssd1 vccd1 vccd1 _16716__1270/HI net1270 sky130_fd_sc_hd__conb_1
XANTENNA__08948__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[25\] vssd1 vssd1 vccd1 vccd1
+ net1407 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ net1119 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XANTENNA_input29_A wbm_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15326__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ net1174 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ net1378 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_13842_ net1083 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
X_16561_ clknet_leaf_29_wb_clk_i net1456 _01434_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13773_ net1135 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XANTENNA__08838__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ _06489_ _06491_ net392 vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15512_ clknet_leaf_121_wb_clk_i _01963_ _00470_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12724_ net977 net979 _04373_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__and4_1
X_16636__1207 vssd1 vssd1 vccd1 vccd1 _16636__1207/HI net1207 sky130_fd_sc_hd__conb_1
X_16492_ clknet_leaf_64_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[27\] _01366_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[27\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15476__CLK clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ clknet_leaf_125_wb_clk_i _01894_ _00401_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12655_ _05793_ _05837_ _05884_ _05931_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12409__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ net259 net2063 net578 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15374_ clknet_leaf_33_wb_clk_i _01825_ _00332_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12586_ net307 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[11\] net475 vssd1
+ vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XANTENNA__09263__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10437__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09802__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14325_ net1120 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ net449 _07125_ _07126_ net429 _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
X_14256_ net1021 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11468_ net442 _07059_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__a21bo_1
X_13207_ team_02_WB.START_ADDR_VAL_REG\[15\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net198 sky130_fd_sc_hd__a21o_1
X_10419_ _06064_ _06071_ net382 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__mux2_1
XANTENNA__12144__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14187_ net1013 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XANTENNA__10176__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _05614_ _06135_ net432 _06016_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13138_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _03131_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_123_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11983__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13764__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ _07434_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12322__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1109 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16497__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07630_ _03482_ _03514_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15819__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ _03443_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16759_ net1313 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_0_18_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09300_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[24\] net870 net834 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09689__A _05337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ net2115 team_02_WB.instance_to_wrap.ramload\[13\] net969 vssd1 vssd1 vccd1
+ vccd1 _02842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _04888_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12319__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09162_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[27\] net669 net659 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[27\]
+ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a221o_1
XANTENNA__09254__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08113_ _03962_ _03994_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13107__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__B1 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09093_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[29\] net770 net758 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13338__C1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ _03889_ _03928_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__xor2_4
Xhold910 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold932 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold943 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10363__A _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12054__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold965 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold976 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold987 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15349__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _05633_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout585_A _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08946_ net898 _04629_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or2_1
XANTENNA__11116__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11116__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] net939 _04328_ _04566_ vssd1
+ vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07828_ _03717_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nand2_1
XANTENNA__10875__B1 team_02_WB.instance_to_wrap.top.aluOut\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15499__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] _03649_ _03647_ _03646_ vssd1
+ vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _06419_ _06420_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__and2_1
XANTENNA__09493__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\] net809 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[21\]
+ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12229__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12440_ net266 net2610 net486 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XANTENNA__09245__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__B2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ net251 net1853 net493 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ net1022 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
X_11322_ _06862_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08442__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15090_ clknet_leaf_11_wb_clk_i _01541_ _00048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14041_ net1062 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
X_11253_ net382 _06761_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _05852_ _05856_ _05858_ _05860_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[3\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_101_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11184_ _06185_ _06189_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13584__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10135_ _05768_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nor2_1
X_15992_ clknet_leaf_126_wb_clk_i _02443_ _00950_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10066_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[6\] net822 net867 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a22o_1
X_14943_ net1009 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XANTENNA__10720__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14874_ net1166 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16613_ clknet_leaf_57_wb_clk_i _02847_ _01486_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ net1143 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ clknet_leaf_6_wb_clk_i net1437 _01417_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13756_ net1097 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
X_10968_ net452 _06143_ _06606_ _06607_ _06608_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11633__C_N team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ _07333_ _07334_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__and2b_2
XFILLER_0_35_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11291__B1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16475_ clknet_leaf_87_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[10\] _01349_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13687_ net1119 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XANTENNA__12139__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10899_ _06142_ _06208_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ clknet_leaf_49_wb_clk_i _01877_ _00384_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12638_ _04826_ _04913_ _04993_ _05156_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__or4_1
XANTENNA__09236__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11978__S net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ clknet_leaf_112_wb_clk_i _01808_ _00315_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_12569_ net250 net2439 net474 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14308_ net1100 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
Xhold206 _02817_ vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15288_ clknet_leaf_123_wb_clk_i _01739_ _00246_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold217 team_02_WB.instance_to_wrap.top.a1.row1\[120\] vssd1 vssd1 vccd1 vccd1 net1615
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _02597_ vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 team_02_WB.START_ADDR_VAL_REG\[23\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net1126 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XANTENNA__16617__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10149__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout708 _04458_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_6
Xfanout719 _04456_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ net165 net951 net902 net1503 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__B _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[12\] net686 net657 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\]
+ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07970__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ net1581 net958 net924 _04522_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08514__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[0\] net715 net710 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07613_ _03501_ _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__and2b_1
X_08593_ net975 _03396_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07544_ _03431_ _03433_ _03434_ _03430_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07475_ team_02_WB.instance_to_wrap.top.a1.instruction\[30\] net1893 net966 vssd1
+ vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
XANTENNA__12049__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout333_A _07035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1075_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[26\] net774 net838 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11888__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09145_ _04824_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout500_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11585__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09076_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] net717 net681 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[29\]
+ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15171__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08027_ _03883_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or2_1
XANTENNA__12723__D team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold740 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold751 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11337__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold762 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold784 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold795 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12512__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[8\] net811 net851 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ _04607_ _04609_ _04611_ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11940_ net258 net2503 net537 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10312__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11871_ net248 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[29\] net545 vssd1
+ vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12748__A _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ net1013 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
X_10822_ net451 _06464_ _06470_ _06458_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14590_ net1200 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09466__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13541_ _03381_ _03382_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10753_ _05929_ net374 _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ clknet_leaf_95_wb_clk_i _02698_ _01217_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input96_A wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08961__A team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ team_02_WB.instance_to_wrap.top.pc\[16\] team_02_WB.instance_to_wrap.top.pc\[15\]
+ _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11798__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15211_ clknet_leaf_20_wb_clk_i _01662_ _00169_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ net328 net2260 net490 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__mux2_1
XANTENNA__11025__B1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13579__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16191_ clknet_leaf_64_wb_clk_i net1609 _01149_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XANTENNA__15514__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15142_ clknet_leaf_13_wb_clk_i _01593_ _00100_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12354_ net301 net2611 net498 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10715__B net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ net424 _06456_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15073_ clknet_leaf_58_wb_clk_i _01524_ _00036_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12285_ net270 net2005 net504 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15664__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14024_ net1097 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ _05658_ _06169_ _06175_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__A _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ net407 _06566_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[5\] net763 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ _06033_ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__or2_1
X_15975_ clknet_leaf_15_wb_clk_i _02426_ _00933_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14926_ net1000 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
X_10049_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[6\] net650 _05708_ vssd1
+ vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a21o_1
XANTENNA__09016__B _04698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11500__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14857_ net1188 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13808_ net1017 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XANTENNA__09457__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14788_ net1176 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11264__B1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16527_ clknet_leaf_29_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[30\]
+ _01401_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ net1013 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ clknet_leaf_57_wb_clk_i net1508 _01332_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15194__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15409_ clknet_leaf_18_wb_clk_i _01860_ _00367_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16389_ clknet_leaf_77_wb_clk_i _02820_ _01263_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.keyCode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11319__A1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07543__D_N team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09901_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[10\] net862 net815 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\]
+ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout505 net507 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_4
Xfanout516 _07213_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08735__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[11\] net731 net699 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[11\]
+ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a221o_1
Xfanout527 _07210_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_8
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_6
XANTENNA__12332__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _07200_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_4
X_09763_ _05423_ _05425_ _05427_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__or4_1
X_08714_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09694_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[14\] net733 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a22o_1
XANTENNA__09696__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09160__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08645_ team_02_WB.instance_to_wrap.top.a1.instruction\[16\] team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ _04439_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout450_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1192_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout548_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ net975 net976 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__and2_1
XANTENNA__09448__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07527_ team_02_WB.instance_to_wrap.top.a1.state\[1\] team_02_WB.instance_to_wrap.top.a1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nor2_2
XANTENNA__12718__D team_02_WB.instance_to_wrap.top.a1.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15537__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout715_A _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14783__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ team_02_WB.instance_to_wrap.top.lcd.currentState\[3\] vssd1 vssd1 vccd1 vccd1
+ _03399_ sky130_fd_sc_hd__inv_2
Xwire906 _04552_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11007__B1 team_02_WB.instance_to_wrap.top.aluOut\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12507__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11558__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[28\] net854 net790 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[28\]
+ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a221o_1
XANTENNA__09620__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09059_ _04722_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ net239 net2013 net524 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold570 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12710__A_N _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ net405 _06116_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__nor2_1
XANTENNA__12242__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13862__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15760_ clknet_leaf_39_wb_clk_i _02211_ _00718_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12972_ _07373_ _07374_ _02865_ net888 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a31o_1
XANTENNA__08956__A team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A wbm_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ net1035 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
Xhold1281 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ net311 net2656 net541 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__10697__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1292 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
X_15691_ clknet_leaf_20_wb_clk_i _02142_ _00649_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ net999 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ net292 net2160 net548 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ net380 _06113_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__nand2_1
X_14573_ net1133 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11785_ net269 net1717 net556 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13524_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[4\]
+ _03368_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__and3_1
X_16312_ clknet_leaf_78_wb_clk_i _02745_ _01255_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10736_ _06385_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16243_ clknet_leaf_93_wb_clk_i _02681_ _01200_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[12\] _03326_ net1175 vssd1
+ vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a21oi_1
X_10667_ _06315_ _06317_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__o21a_1
XANTENNA__12417__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10726__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12406_ net258 net1985 net489 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16174_ clknet_leaf_66_wb_clk_i _02620_ _01132_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ team_02_WB.instance_to_wrap.top.a1.row1\[109\] _03273_ _03285_ team_02_WB.instance_to_wrap.top.a1.row1\[101\]
+ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10598_ team_02_WB.instance_to_wrap.top.pc\[21\] _06248_ vssd1 vssd1 vccd1 vccd1
+ _06250_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15125_ clknet_leaf_123_wb_clk_i _01576_ _00083_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12337_ net248 net1704 net497 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ clknet_leaf_91_wb_clk_i _01507_ _00019_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12268_ _04576_ _07188_ _07194_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or3_1
XANTENNA__12660__B _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ net1114 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11219_ _06027_ _06841_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12152__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12199_ net358 net2341 net516 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09390__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10180__B _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15958_ clknet_leaf_108_wb_clk_i _02409_ _00916_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09678__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11485__B1 _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14909_ net1146 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15889_ clknet_leaf_19_wb_clk_i _02340_ _00847_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08430_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\] net917 vssd1 vssd1 vccd1
+ vccd1 _04293_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08361_ _04231_ _04233_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12985__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _04133_ _04137_ _04169_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__and3_1
XANTENNA__09850__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12327__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09602__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _06956_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12062__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1205_A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 _07055_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
Xfanout346 net349 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input3_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 _07135_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
X_09815_ net607 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[12\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__09381__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout368 net371 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_4
Xfanout379 net381 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
XANTENNA_fanout665_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\] net648 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[13\]
+ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a221o_1
XANTENNA__09669__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[15\] net841 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[15\]
+ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08628_ net931 net740 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08559_ net83 net1624 net892 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12976__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11570_ net454 _06155_ _07160_ _04604_ _07162_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a221o_1
XANTENNA__09841__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ _05591_ _05613_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12237__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14018__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ team_02_WB.instance_to_wrap.ramload\[13\] net983 vssd1 vssd1 vccd1 vccd1
+ team_02_WB.instance_to_wrap.top.ru.dmmload_co\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_33_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ _05768_ net369 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand2_1
XANTENNA__08016__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ _03154_ _03156_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or3_1
XANTENNA__13857__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ _06033_ _06035_ _05114_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o21a_1
XANTENNA__12761__A _05175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12122_ net302 net2296 net588 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input59_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08450__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12053_ net269 net2315 net528 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10506__A2 _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ team_02_WB.instance_to_wrap.top.pc\[24\] _06341_ vssd1 vssd1 vccd1 vccd1
+ _06642_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09372__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15702__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 _04667_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_8
X_15812_ clknet_leaf_19_wb_clk_i _02263_ _00770_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout891 net894 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_4
X_16792_ net1346 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
XANTENNA__07590__A team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ _02870_ _02986_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__xnor2_1
X_15743_ clknet_leaf_26_wb_clk_i _02194_ _00701_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ net255 net2272 net542 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15674_ clknet_leaf_120_wb_clk_i _02125_ _00632_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12886_ _02918_ _02919_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14625_ net1157 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
X_11837_ net243 net1818 net550 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14556_ net1098 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
X_11768_ _04577_ _07190_ _07194_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__or3_4
XANTENNA__09832__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13507_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[8\] _03358_
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[10\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16208__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _04722_ net371 vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ net1111 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__A _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ net360 net1852 net570 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16226_ clknet_leaf_29_wb_clk_i _02671_ _01183_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13438_ _03303_ _03307_ _03317_ net1176 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_113_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08399__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11986__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16157_ clknet_leaf_7_wb_clk_i net1554 _01115_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13369_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] _03271_ vssd1 vssd1 vccd1
+ vccd1 _03272_ sky130_fd_sc_hd__nand2_1
XANTENNA__16358__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15232__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15108_ clknet_leaf_55_wb_clk_i _01559_ _00066_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16088_ clknet_leaf_80_wb_clk_i _02534_ _01046_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07930_ _03762_ _03807_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__xor2_1
X_15039_ net1154 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09899__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09363__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _03746_ _03747_ _03749_ _03744_ _03707_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] net824 net860 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07792_ net341 _03679_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] vssd1 vssd1
+ vccd1 vccd1 _03683_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09531_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[18\] net689 net641 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a22o_1
XANTENNA__09115__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09462_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] net785 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10130__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08874__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04270_ _04276_ net991 vssd1
+ vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[22\] net851 net779 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[22\]
+ _05054_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout246_A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ _04185_ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08535__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12057__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ _04146_ _04148_ _04152_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout413_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1155_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10085__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11896__S net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13677__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout782_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15725__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1108 net1113 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_4
Xfanout1119 net1122 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_4
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09354__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15875__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ _05390_ _05392_ _05394_ _05396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[14\]
+ sky130_fd_sc_hd__or4_4
XFILLER_0_9_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ team_02_WB.instance_to_wrap.top.i_ready net988 vssd1 vssd1 vccd1 vccd1 _07364_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10121__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12671_ _06963_ _06966_ _06986_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12756__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__B1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ net1037 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
X_11622_ net312 net2371 net577 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15390_ clknet_leaf_3_wb_clk_i _01841_ _00348_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11621__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ net1087 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11553_ net440 _07144_ _07145_ net426 _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ net366 _05975_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15255__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14272_ net1079 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
X_11484_ _06714_ _07083_ net409 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__mux2_1
X_16011_ clknet_leaf_20_wb_clk_i _02462_ _00969_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13223_ team_02_WB.START_ADDR_VAL_REG\[31\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net216 sky130_fd_sc_hd__a21o_1
XFILLER_0_122_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12716__A3 _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _05378_ net372 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nand2_1
Xwire599 _05743_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10188__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09593__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ _03398_ net895 _03145_ net1183 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a211o_2
XFILLER_0_27_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10366_ _05572_ _06018_ _05570_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a21o_1
XANTENNA__10723__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ net248 net2657 net587 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
X_13085_ _07405_ _07428_ _07429_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10297_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[1\] net845 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12036_ net594 _07190_ _07205_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__or3_1
XANTENNA__09345__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11152__A2 team_02_WB.instance_to_wrap.top.aluOut\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12430__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775_ net1329 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13987_ net1068 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15726_ clknet_leaf_42_wb_clk_i _02177_ _00684_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12938_ _02878_ _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__and2_1
XANTENNA__08856__B2 team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15657_ clknet_leaf_31_wb_clk_i _02108_ _00615_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16030__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ team_02_WB.instance_to_wrap.top.pc\[16\] _06266_ vssd1 vssd1 vccd1 vccd1
+ _02903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14608_ net1196 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
X_15588_ clknet_leaf_55_wb_clk_i _02039_ _00546_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14539_ net1026 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XANTENNA__14881__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10966__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] _03869_ _03903_ vssd1 vssd1
+ vccd1 vccd1 _03948_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15748__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16209_ clknet_leaf_28_wb_clk_i _02654_ _01166_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09584__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16809__1363 vssd1 vssd1 vccd1 vccd1 _16809__1363/HI net1363 sky130_fd_sc_hd__conb_1
XANTENNA__08792__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ net883 _04639_ _04641_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_4
XFILLER_0_122_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07913_ _03801_ _03803_ _03797_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_2
XANTENNA__15898__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ team_02_WB.instance_to_wrap.top.a1.instruction\[8\] team_02_WB.instance_to_wrap.top.a1.instruction\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07844_ _03702_ _03716_ _03734_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12340__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10550__A_N _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15128__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _03662_ _03664_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__xor2_1
X_09514_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] net819 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10103__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[20\] net724 net660 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\]
+ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout628_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15278__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _05042_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nor2_4
XFILLER_0_69_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08327_ _04202_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14791__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08258_ _04114_ _04116_ _04136_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout997_A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ _04066_ _04068_ _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3_1
XANTENNA__12515__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10220_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[3\] net727 net663 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\]
+ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a221o_1
XANTENNA__09575__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08783__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10151_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\] net814 net797 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\]
+ _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09327__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[6\] net803 net799 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\]
+ _05727_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a221o_1
X_13910_ net1109 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XANTENNA__12250__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1175 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ net1029 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XANTENNA__16053__CLK clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ clknet_leaf_39_wb_clk_i net1459 _01433_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13772_ net1003 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13292__C1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ net383 _06487_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__nand2_1
XANTENNA__08964__A team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15511_ clknet_leaf_119_wb_clk_i _01962_ _00469_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12723_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] team_02_WB.instance_to_wrap.top.a1.instruction\[30\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] team_02_WB.instance_to_wrap.top.a1.instruction\[28\]
+ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__and4_1
X_16491_ clknet_leaf_58_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[26\] _01365_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[26\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _05838_ _05933_ _07273_ _07281_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__or4b_1
X_15442_ clknet_leaf_25_wb_clk_i _01893_ _00400_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ net256 net2238 net579 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15373_ clknet_leaf_24_wb_clk_i _01824_ _00331_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ net299 net2546 net473 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14324_ net1039 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ _06006_ net454 net446 _06003_ _07129_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ net1124 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12425__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11467_ net434 _07065_ _07066_ net448 _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10734__A _05503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ team_02_WB.START_ADDR_VAL_REG\[14\] _04356_ vssd1 vssd1 vccd1 vccd1 net197
+ sky130_fd_sc_hd__and2_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ _06067_ _06070_ net364 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__mux2_1
X_14186_ net1036 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
X_11398_ net422 _06596_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__nor2_1
X_13137_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[1\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10349_ _05930_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_1
XANTENNA__09318__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ _07399_ _07400_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__nand2_1
X_12019_ net324 net2267 net468 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12160__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10333__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14876__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _03447_ _03450_ _03449_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13283__C1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16758_ net1312 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_57_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15420__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16546__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15709_ clknet_leaf_113_wb_clk_i _02160_ _00667_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_07491_ net974 team_02_WB.instance_to_wrap.ramload\[14\] net969 vssd1 vssd1 vccd1
+ vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XANTENNA__09689__B _05355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07501__A1 team_02_WB.instance_to_wrap.ramload\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16689_ net1243 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_14_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ net898 _04908_ _04630_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] net725 net645 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _03993_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09092_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[29\] net810 net782 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[29\]
+ _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13338__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ _03910_ _03926_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a21o_2
XFILLER_0_71_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12335__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09557__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold944 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold955 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold977 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09994_ _05636_ net603 net899 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__mux2_1
Xhold988 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09309__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ net898 _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_2
XANTENNA__16076__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] net915 _04312_ net959 vssd1
+ vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _03702_ _03709_ _03710_ _03715_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__or4bb_2
XANTENNA__10875__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14786__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07758_ _03408_ net350 vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ _03573_ _03579_ _03574_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10819__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15913__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] net853 net769 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[22\] net718 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[22\]
+ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12370_ net249 net2456 net493 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ _05484_ _06861_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ net1056 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net387 _06872_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10203_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[3\] net824 net796 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\]
+ _05859_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a221o_1
XANTENNA__16419__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11183_ _06185_ _06807_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11569__A2_N _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10134_ net899 net597 _05772_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a21o_1
X_15991_ clknet_leaf_116_wb_clk_i _02442_ _00949_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] net749 _05724_ vssd1
+ vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__o21a_2
X_14942_ net1007 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XANTENNA__10315__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15443__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16569__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ net1188 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16612_ clknet_leaf_61_wb_clk_i _02846_ _01485_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ net1082 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10618__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16543_ clknet_leaf_0_wb_clk_i net1455 _01416_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ net1046 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XANTENNA__15593__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ net448 _06603_ _06597_ net439 vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a2bb2o_1
X_16808__1362 vssd1 vssd1 vccd1 vccd1 _16808__1362/HI net1362 sky130_fd_sc_hd__conb_1
XFILLER_0_85_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07495__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12647__C _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _07328_ _07327_ team_02_WB.instance_to_wrap.top.aluOut\[31\] vssd1 vssd1
+ vccd1 vccd1 _07334_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16474_ clknet_leaf_91_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[9\] _01348_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[9\] sky130_fd_sc_hd__dfrtp_1
X_13686_ net1111 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
X_10898_ net439 _06532_ _06538_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15425_ clknet_leaf_0_wb_clk_i _01876_ _00383_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _05934_ _06006_ _06011_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15356_ clknet_leaf_48_wb_clk_i _01807_ _00314_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12568_ net246 net2673 net474 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09787__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14307_ net1069 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
X_11519_ net345 net1804 net584 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12155__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ team_02_WB.instance_to_wrap.top.a1.instruction\[7\] net594 _07187_ _07204_
+ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__and4_4
X_15287_ clknet_leaf_118_wb_clk_i _01738_ _00245_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold207 net150 vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold218 team_02_WB.instance_to_wrap.top.a1.row1\[10\] vssd1 vssd1 vccd1 vccd1 net1616
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold229 team_02_WB.instance_to_wrap.top.a1.row1\[123\] vssd1 vssd1 vccd1 vccd1 net1627
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ net1021 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11994__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14169_ net1064 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout709 _04458_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[27\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[27\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
XANTENNA__07970__B2 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11503__C1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08661_ net747 _04449_ _04455_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__and3_4
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07612_ _03460_ _03502_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15936__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08592_ net973 net975 _03396_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07543_ team_02_WB.instance_to_wrap.top.a1.dataIn\[23\] team_02_WB.instance_to_wrap.top.a1.dataIn\[21\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[20\] team_02_WB.instance_to_wrap.top.a1.dataIn\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10639__A team_02_WB.instance_to_wrap.top.pc\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07474_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] team_02_WB.instance_to_wrap.ramload\[31\]
+ net965 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[26\] net871 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\]
+ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12854__A team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09144_ _04804_ _04823_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09778__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15316__CLK clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09075_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\] net725 net658 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a22o_1
XANTENNA__12065__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08026_ _03846_ _03878_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold730 team_02_WB.instance_to_wrap.top.a1.row2\[25\] vssd1 vssd1 vccd1 vccd1 net2128
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout695_A _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold763 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold774 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15466__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[8\] net871 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ _05637_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout862_A _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08928_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[31\] net720 net712 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\]
+ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09702__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08859_ team_02_WB.instance_to_wrap.top.edg2.flip2 _04283_ team_02_WB.instance_to_wrap.top.edg2.flip1
+ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nor3b_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ net242 net2545 net545 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ _04785_ net453 _06468_ net436 _06469_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07477__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13540_ net2062 _03379_ net884 vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10752_ _05975_ net374 vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13471_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[0\] net873 vssd1 vssd1 vccd1
+ vccd1 _02786_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ team_02_WB.instance_to_wrap.top.pc\[14\] _06334_ vssd1 vssd1 vccd1 vccd1
+ _06335_ sky130_fd_sc_hd__and2_1
XANTENNA__12764__A _05247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15210_ clknet_leaf_51_wb_clk_i _01661_ _00168_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12422_ net311 net2470 net490 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__mux2_1
XANTENNA__11025__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ clknet_leaf_63_wb_clk_i _02636_ _01148_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input89_A wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15141_ clknet_leaf_127_wb_clk_i _01592_ _00099_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12353_ net292 net2200 net496 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ net413 _06463_ _06919_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__o21ba_1
X_15072_ clknet_leaf_57_wb_clk_i _01523_ _00035_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[25\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_26_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12284_ net325 net2009 net504 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08729__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ net1152 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11235_ net324 net2428 net582 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10000__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _06792_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__inv_2
XANTENNA__09941__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10117_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[5\] net791 net776 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\]
+ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a221o_1
X_15974_ clknet_leaf_3_wb_clk_i _02425_ _00932_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11097_ _05156_ _06032_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10048_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[6\] net666 net630 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a22o_1
X_14925_ net1001 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[10\] vssd1 vssd1 vccd1 vccd1
+ net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14856_ net1191 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ net1129 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10459__A _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14787_ net1184 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
X_11999_ net1752 _07153_ net532 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
X_16526_ clknet_leaf_39_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[29\]
+ _01400_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10067__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13738_ net1036 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16457_ clknet_leaf_64_wb_clk_i net1497 _01331_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13669_ net1089 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ clknet_leaf_39_wb_clk_i _01859_ _00366_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_16388_ clknet_leaf_73_wb_clk_i _02819_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15339_ clknet_leaf_16_wb_clk_i _01790_ _00297_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[10\] net795 net775 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10922__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09393__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[11\] net718 net631 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a22o_1
Xfanout517 _07213_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_4
XANTENNA__09932__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout528 net531 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_8
Xfanout539 _07203_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\] net861 net789 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[13\]
+ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a221o_1
X_08713_ net750 _04509_ _04508_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o21a_4
X_09693_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] net729 net721 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[14\]
+ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08644_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04439_ vssd1 vssd1
+ vccd1 vccd1 _04441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16114__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__inv_2
XANTENNA__10369__A _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_A _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1185_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] net990 _03417_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand4b_2
XANTENNA__10058__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09999__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11899__S net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ team_02_WB.instance_to_wrap.top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1
+ _03398_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout708_A _04458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11007__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11558__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08959__B1 _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] net870 net846 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ net901 team_02_WB.instance_to_wrap.top.DUT.read_data2\[30\] net593 vssd1
+ vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08009_ _03870_ _03871_ net241 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21oi_2
Xhold560 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12523__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
X_16807__1361 vssd1 vssd1 vccd1 vccd1 _16807__1361/HI net1361 sky130_fd_sc_hd__conb_1
X_11020_ _06040_ net452 _06655_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a211o_1
XANTENNA__09384__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold593 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09923__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09136__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ _02967_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09687__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12759__A _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1260 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08956__B team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ net1033 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
Xhold1271 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ net308 net2023 net543 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
Xhold1282 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11494__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1293 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ clknet_leaf_45_wb_clk_i _02141_ _00648_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ net1008 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ net285 net2627 net550 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XANTENNA__13092__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _06106_ _06110_ net365 vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ net1005 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
X_11784_ net325 net2159 net556 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16311_ clknet_leaf_77_wb_clk_i _02744_ _01254_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_13523_ net1614 _03368_ _03370_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10735_ _05461_ net369 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__nand2_1
XANTENNA__08662__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11602__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16242_ clknet_leaf_93_wb_clk_i _02680_ _01199_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_10666_ _06315_ _06317_ _04416_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__a21oi_1
X_13454_ _03326_ _03327_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nor2_1
XANTENNA__10726__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12405_ net254 net2219 net489 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16173_ clknet_leaf_66_wb_clk_i _02619_ _01131_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
X_13385_ team_02_WB.instance_to_wrap.top.a1.row1\[13\] _03217_ _03221_ _03226_ team_02_WB.instance_to_wrap.top.a1.row1\[61\]
+ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10597_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__inv_2
XANTENNA__10221__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15124_ clknet_leaf_53_wb_clk_i _01575_ _00082_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12336_ net244 net1954 net497 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15055_ clknet_leaf_89_wb_clk_i _01506_ _00018_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_12267_ net236 net2414 net511 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10742__A _05677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11218_ _05318_ _06026_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__nor2_1
X_14006_ net1109 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XANTENNA__09914__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ net351 net2668 net516 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ net912 _06776_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16137__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15957_ clknet_leaf_115_wb_clk_i _02408_ _00915_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12669__A _07005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ net1147 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__10288__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15888_ clknet_leaf_39_wb_clk_i _02339_ _00846_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14839_ net1169 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08360_ _04227_ _04229_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12985__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16509_ clknet_leaf_1_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[12\]
+ _01383_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_08291_ _04137_ _04169_ _04133_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_131_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12201__A3 team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12343__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout303 _06780_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout314 _06996_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_1
Xfanout325 _06856_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
XANTENNA_fanout393_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _07055_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
X_09814_ _05473_ _05477_ _05478_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nor4_2
Xfanout347 net349 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout358 net361 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1100_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[13\] net628 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout560_A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15504__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09676_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] net861 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08627_ _04360_ _04421_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14794__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08558_ net94 net1693 net893 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15654__CLK clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07509_ net2631 net119 _00011_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12518__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08489_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _04276_ vssd1 vssd1 vccd1
+ vccd1 _04326_ sky130_fd_sc_hd__nor2_2
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10520_ _05544_ _05569_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10451_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10203__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13170_ _03144_ _03146_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11400__A1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ _05154_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ net291 net1864 net586 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12253__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ net324 net2039 net528 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold390 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _06243_ _06303_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_73_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout870 _04642_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_4
X_15811_ clknet_leaf_43_wb_clk_i _02262_ _00769_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout881 _04667_ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ net1345 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XANTENNA__15184__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout892 net894 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15742_ clknet_leaf_4_wb_clk_i _02193_ _00700_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12954_ _07368_ _07369_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11467__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1090 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10675__C1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ net253 net2281 net542 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
X_15673_ clknet_leaf_107_wb_clk_i _02124_ _00631_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12885_ team_02_WB.instance_to_wrap.top.pc\[7\] _05725_ vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_16_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14624_ net1157 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
X_11836_ net238 net2284 net550 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14555_ net1060 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XANTENNA__12428__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ net234 net2654 net561 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XANTENNA__10978__B1 team_02_WB.instance_to_wrap.top.aluOut\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13506_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[5\] team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[6\]
+ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[7\] vssd1 vssd1 vccd1
+ vccd1 _03358_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10718_ net378 _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__nor2_1
X_14486_ net1108 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11698_ net353 net1921 net568 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16225_ clknet_leaf_7_wb_clk_i _02670_ _01182_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13437_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\] _03301_ net1587 vssd1 vssd1
+ vccd1 vccd1 _03317_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ _06250_ _06300_ _06247_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09596__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16156_ clknet_leaf_7_wb_clk_i net1561 _01114_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13368_ net985 _03215_ _03211_ team_02_WB.instance_to_wrap.top.lcd.nextState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_24_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15107_ clknet_leaf_43_wb_clk_i _01558_ _00065_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12163__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net285 net2286 net500 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
XANTENNA__10472__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16087_ clknet_leaf_79_wb_clk_i _02533_ _01045_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13299_ _03146_ _03155_ _02780_ _03170_ _03148_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__o311a_1
XFILLER_0_126_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09348__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15038_ net1154 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15527__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _03707_ _03749_ _03748_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07791_ _03648_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09530_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[18\] net658 _05201_ vssd1
+ vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09461_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08412_ team_02_WB.instance_to_wrap.top.a1.state\[0\] _04268_ vssd1 vssd1 vccd1 vccd1
+ _04279_ sky130_fd_sc_hd__and2_2
X_09392_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[22\] net880 _05065_ _05067_
+ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16806__1360 vssd1 vssd1 vccd1 vccd1 _16806__1360/HI net1360 sky130_fd_sc_hd__conb_1
XFILLER_0_30_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08343_ _04208_ _04215_ _04202_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12338__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14119__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11091__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04153_ vssd1 vssd1 vccd1
+ vccd1 _04154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13958__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09587__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08551__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11478__A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13135__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09339__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1109 net1113 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout942_A _07365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ _03841_ _03860_ _03842_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09728_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[14\] net758 net754 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[14\]
+ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a221o_1
XANTENNA__12102__A team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[15\] net701 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12670_ _07025_ _07043_ _07296_ _07297_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__or4b_1
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11621_ net307 net2479 net579 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13071__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12248__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14029__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14340_ net1146 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
X_11552_ _05934_ net454 _06135_ _05932_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09290__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16695__1249 vssd1 vssd1 vccd1 vccd1 _16695__1249/HI net1249 sky130_fd_sc_hd__conb_1
X_10503_ _06112_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ net1112 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
X_11483_ _06715_ _07083_ net409 vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16010_ clknet_leaf_45_wb_clk_i _02461_ _00968_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09578__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input71_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ team_02_WB.START_ADDR_VAL_REG\[30\] net997 net933 vssd1 vssd1 vccd1 vccd1
+ net215 sky130_fd_sc_hd__a21o_1
X_10434_ _05337_ net367 vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nand2_1
XANTENNA__09042__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11385__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ team_02_WB.instance_to_wrap.top.lcd.currentState\[4\] net895 vssd1 vssd1
+ vccd1 vccd1 _03145_ sky130_fd_sc_hd__nor2_1
X_10365_ _06015_ _06017_ _05614_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ net243 net1958 net587 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
X_13084_ _07366_ _03095_ team_02_WB.instance_to_wrap.top.pc\[9\] net945 vssd1 vssd1
+ vccd1 vccd1 _01507_ sky130_fd_sc_hd__a2bb2o_1
X_10296_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] net793 _05948_ _05950_
+ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a211o_1
X_12035_ net235 net2695 net469 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09750__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11327__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16774_ net1328 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
X_13986_ net1088 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
X_15725_ clknet_leaf_24_wb_clk_i _02176_ _00683_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12937_ _02879_ _02970_ _02880_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10112__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08856__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15656_ clknet_leaf_56_wb_clk_i _02107_ _00614_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12868_ team_02_WB.instance_to_wrap.top.pc\[17\] _06263_ vssd1 vssd1 vccd1 vccd1
+ _02902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14607_ net1196 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
X_11819_ net285 net2233 net553 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
X_15587_ clknet_leaf_43_wb_clk_i _02038_ _00545_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12158__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__A _04602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13062__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ _05725_ _05722_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14538_ net1051 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XANTENNA__16325__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11997__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14469_ net1089 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
XANTENNA__12682__A _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09569__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ clknet_leaf_37_wb_clk_i _02653_ _01165_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09033__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ clknet_leaf_129_wb_clk_i net1529 _01097_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ team_02_WB.instance_to_wrap.top.a1.instruction\[20\] net883 _04635_ _04644_
+ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07912_ _03774_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08892_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04429_ vssd1 vssd1
+ vccd1 vccd1 _04577_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07843_ _03701_ _03733_ _03692_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a21o_1
XANTENNA__13018__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _03631_ _03636_ _03662_ net350 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__or4b_1
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09513_ _05179_ _05181_ _05183_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__or4_1
XANTENNA__11834__C_N team_02_WB.instance_to_wrap.top.a1.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08847__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1098_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\] net656 net628 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09231__A _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _05044_ _05046_ _05048_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__or4_2
XANTENNA__12068__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A _07212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11064__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ _04187_ _04194_ _04196_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08257_ _04134_ _04126_ _04123_ _04129_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__and4b_1
XANTENNA__08480__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11700__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08188_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] _04071_ vssd1 vssd1 vccd1
+ vccd1 _04072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09024__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout892_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13200__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08783__B2 _04548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[4\] net861 net853 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[6\] net819 net779 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ _05726_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a221o_1
XANTENNA__12531__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net1016 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ net1013 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XANTENNA__08838__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _06484_ _06488_ net390 vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15510_ clknet_leaf_112_wb_clk_i _01961_ _00468_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ net972 _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16490_ clknet_leaf_57_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[25\] _01364_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[25\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09141__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ clknet_leaf_17_wb_clk_i _01892_ _00399_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12653_ _05571_ _05614_ _05657_ net425 vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ net250 net2474 net578 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09799__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ clknet_leaf_52_wb_clk_i _01823_ _00330_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12584_ net293 net1770 net472 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__mux2_1
XANTENNA__09263__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15372__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14323_ net1102 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
X_11535_ net412 net438 _06756_ net432 _05884_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__a32o_1
XANTENNA__16498__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12706__S team_02_WB.instance_to_wrap.top.aluOut\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11610__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14254_ net1065 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
X_11466_ net423 net437 _06687_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13205_ team_02_WB.START_ADDR_VAL_REG\[13\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net196 sky130_fd_sc_hd__a21o_1
XFILLER_0_106_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10417_ _06068_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11397_ net413 _06602_ _07004_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__o21ba_1
X_14185_ net1011 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XANTENNA__10030__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _04343_ _04551_ team_02_WB.instance_to_wrap.wb.curr_state\[2\] _03404_ vssd1
+ vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_123_1654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10348_ _05931_ _05932_ _05976_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12441__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _05931_ _05932_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__nor2_1
X_13067_ _06972_ net227 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nor2_1
XANTENNA__09723__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ net320 net2712 net471 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ net152 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ net1311 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
XANTENNA__08829__A2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ net1031 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XANTENNA__11581__A _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ clknet_leaf_62_wb_clk_i _02159_ _00666_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_07490_ team_02_WB.instance_to_wrap.top.a1.instruction\[15\] net1647 net970 vssd1
+ vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__mux2_1
XANTENNA__08227__D_N team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16688_ net1242 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_53_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15639_ clknet_leaf_118_wb_clk_i _02090_ _00597_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15715__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14892__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09160_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[27\] net737 net729 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[27\]
+ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09254__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ _03920_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\] net778 net767 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ _03929_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09006__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold912 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold934 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold945 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10021__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__B2 _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold967 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09962__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold978 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net601 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[8\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net749 _04628_ vssd1
+ vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o21a_2
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12351__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09714__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net1552 _04565_ net825 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _07226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16694__1248 vssd1 vssd1 vccd1 vccd1 _16694__1248/HI net1248 sky130_fd_sc_hd__conb_1
X_07826_ _03692_ _03701_ _03709_ _03690_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a31oi_4
XANTENNA__15245__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07757_ _03646_ _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout640_A _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout738_A _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07688_ _03530_ _03557_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09493__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15395__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\] net785 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[21\]
+ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\] net708 net678 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__a22o_1
XANTENNA__09245__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ _04153_ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09289_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[24\] net725 net717 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11430__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ net291 net2397 net582 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11251_ _06815_ _06871_ net376 vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10012__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10202_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[3\] net868 net877 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a22o_1
XANTENNA__09953__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11182_ _05316_ _06027_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ net899 net597 _05772_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12261__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15990_ clknet_leaf_109_wb_clk_i _02441_ _00948_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09705__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A wbm_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ net462 _05679_ _05723_ net456 net740 vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a221o_1
X_14941_ net1007 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
X_14872_ net1190 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ clknet_leaf_60_wb_clk_i _02845_ _01484_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13823_ net1125 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15738__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11605__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ clknet_leaf_37_wb_clk_i net1439 _01415_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13754_ net1038 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
X_10966_ _06043_ net430 net445 _04952_ _06583_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__a221o_1
XANTENNA__09484__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12705_ _07323_ _07324_ _07322_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16473_ clknet_leaf_88_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[8\] _01347_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[8\] sky130_fd_sc_hd__dfrtp_1
X_13685_ net1120 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _04869_ net430 net445 _04867_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15424_ clknet_leaf_9_wb_clk_i _01875_ _00382_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ _06987_ _07007_ _07027_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__or4_1
XANTENNA__15888__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ clknet_leaf_104_wb_clk_i _01806_ _00313_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12436__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ net242 net2608 net474 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ net1088 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ _04583_ team_02_WB.instance_to_wrap.top.aluOut\[4\] _07115_ vssd1 vssd1 vccd1
+ vccd1 _07116_ sky130_fd_sc_hd__a21o_4
XFILLER_0_103_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15286_ clknet_leaf_110_wb_clk_i _01737_ _00244_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ net234 net1952 net483 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__mux2_1
Xhold208 team_02_WB.START_ADDR_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15118__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold219 net125 vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ net1030 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ net914 _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12960__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__B2 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ net1055 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ net231 _03123_ _07413_ _03121_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12171__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10480__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ net1148 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XANTENNA__15268__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14887__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ net746 _04442_ _04455_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__and3_4
XFILLER_0_59_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] _03465_ _03472_ _03455_ vssd1
+ vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__or4b_1
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16809_ net1363 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08591_ _04364_ _04368_ net887 _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07542_ team_02_WB.instance_to_wrap.top.a1.dataIn\[31\] team_02_WB.instance_to_wrap.top.a1.dataIn\[30\]
+ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09475__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ team_02_WB.instance_to_wrap.top.ru.dmmWen net984 vssd1 vssd1 vccd1 vccd1
+ _03413_ sky130_fd_sc_hd__nor2_1
XANTENNA__07486__A1 team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09212_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\] net847 net768 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12854__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ _04804_ _04823_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09074_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\] net689 net684 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[29\]
+ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08025_ _03875_ _03877_ _03880_ net241 vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold720 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold731 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold753 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold764 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold775 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _04468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12081__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[8\] net819 net835 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08927_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[31\] net688 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout855_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net7 net948 net922 net1686 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07809_ _03666_ _03696_ _03698_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__or3_1
X_08789_ net1620 net953 net904 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[31\]
+ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10820_ _04783_ net430 net445 _04784_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09466__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _06399_ _06401_ net366 vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_98_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _03137_ _03309_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08734__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10682_ team_02_WB.instance_to_wrap.top.pc\[13\] team_02_WB.instance_to_wrap.top.pc\[12\]
+ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__and3_1
XANTENNA__12764__B _05256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net308 net2574 net491 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12256__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15140_ clknet_leaf_19_wb_clk_i _01591_ _00098_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12352_ net285 net2314 net497 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ net420 _06467_ _06919_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15071_ clknet_leaf_57_wb_clk_i _01522_ _00034_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[24\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net320 net2693 net506 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09926__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022_ net1139 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
X_11234_ net461 team_02_WB.instance_to_wrap.top.aluOut\[16\] _06840_ vssd1 vssd1 vccd1
+ vccd1 _06856_ sky130_fd_sc_hd__o21a_4
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11165_ net395 _06791_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10116_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[5\] net795 net771 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a22o_1
X_15973_ clknet_leaf_127_wb_clk_i _02424_ _00931_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11096_ net289 net2188 net582 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[6\] net682 net673 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[6\]
+ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a221o_1
X_14924_ net1001 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold80 _02584_ vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[2\] vssd1 vssd1 vccd1 vccd1
+ net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_14855_ net1161 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13806_ net1064 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14786_ net1180 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11998_ net1914 net356 net535 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XANTENNA__09457__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16525_ clknet_leaf_29_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[28\]
+ _01399_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13737_ net1011 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10949_ _06444_ _06450_ net387 vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16456_ clknet_leaf_64_wb_clk_i net1518 _01330_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13668_ net1101 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ clknet_leaf_33_wb_clk_i _01858_ _00365_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12619_ _06677_ _06773_ _07246_ _06937_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__or4b_1
X_16387_ clknet_leaf_73_wb_clk_i _02818_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12166__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ net1118 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10224__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08968__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15338_ clknet_leaf_45_wb_clk_i _01789_ _00296_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09090__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16693__1247 vssd1 vssd1 vccd1 vccd1 _16693__1247/HI net1247 sky130_fd_sc_hd__conb_1
XFILLER_0_129_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15269_ clknet_leaf_126_wb_clk_i _01720_ _00227_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09917__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout507 _07217_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_8
X_09830_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[11\] net739 net654 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\]
+ _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout518 _07213_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_8
Xfanout529 net531 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_4
XFILLER_0_123_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09761_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] net805 net829 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a22o_1
X_08712_ team_02_WB.instance_to_wrap.top.a1.instruction\[21\] net615 _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a22o_2
X_09692_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[14\] net674 net665 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09696__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] _04439_ vssd1 vssd1
+ vccd1 vccd1 _04440_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout269_A _06891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ net977 net979 _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__or3_2
XFILLER_0_89_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09448__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10369__B _05440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07525_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] net990 _03417_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12865__A team_02_WB.instance_to_wrap.top.pc\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout436_A _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1178_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07456_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1
+ _03397_ sky130_fd_sc_hd__inv_2
XANTENNA__08554__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12076__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10385__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08959__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10215__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[28\] net823 net778 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a22o_1
XANTENNA__15433__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16559__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ _04726_ _04735_ _04738_ _04740_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[30\]
+ sky130_fd_sc_hd__or4_4
X_08008_ _03895_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__or2_1
Xhold550 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A team_02_WB.instance_to_wrap.top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] vssd1 vssd1 vccd1 vccd1
+ net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold583 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold594 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold383_A team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09959_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[8\] net693 net657 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a22o_1
X_12970_ _02884_ _02885_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__nand2_1
Xhold1250 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09687__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1261 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11921_ net300 net1994 net540 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
Xhold1272 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net2681
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
X_14640_ net1007 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
X_11852_ net267 net1931 net548 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10803_ _06450_ _06451_ net387 vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10994__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14571_ net1014 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
X_11783_ net320 net2336 net559 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12775__A _05493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16310_ clknet_leaf_78_wb_clk_i _02743_ _01253_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13522_ net1614 _03368_ net885 vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10734_ _05503_ net374 vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ clknet_leaf_79_wb_clk_i _02679_ _01198_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13453_ net1652 _03325_ net994 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o21ai_1
X_10665_ team_02_WB.instance_to_wrap.top.pc\[31\] _06316_ vssd1 vssd1 vccd1 vccd1
+ _06317_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14990__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ net252 net1947 net489 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__mux2_1
X_16172_ clknet_leaf_66_wb_clk_i _02618_ _01130_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09072__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13384_ team_02_WB.instance_to_wrap.top.lcd.nextState\[5\] _03398_ _03225_ _03272_
+ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_84_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10596_ net928 _04509_ net590 vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__a21o_2
XANTENNA__09611__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15123_ clknet_leaf_126_wb_clk_i _01574_ _00081_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12335_ net237 net1940 net496 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__mux2_1
XANTENNA__15926__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15054_ clknet_leaf_89_wb_clk_i _01505_ _00017_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_12266_ net361 net2473 net508 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
XANTENNA__10509__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10742__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ net1118 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12660__D _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _06263_ net743 _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12197_ net355 net2184 net519 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
X_11148_ _06338_ _06775_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15956_ clknet_leaf_47_wb_clk_i _02407_ _00914_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12131__A0 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ net400 _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__or2_1
XANTENNA__09678__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net1188 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
X_15887_ clknet_leaf_33_wb_clk_i _02338_ _00845_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ net1170 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14769_ net1179 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XANTENNA__12685__A _06569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16508_ clknet_leaf_37_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[11\]
+ _01382_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12985__A2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15456__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ _04159_ _04167_ _04144_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09850__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ clknet_leaf_89_wb_clk_i net1565 _01313_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09063__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09602__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08810__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 _06780_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_1
XFILLER_0_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout315 net318 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
Xfanout326 net329 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_2
Xfanout337 net340 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
X_09813_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[12\] net791 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[12\]
+ _05464_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a221o_1
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
Xfanout359 net361 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09744_ _05404_ _05406_ _05408_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__or4_2
XANTENNA__09669__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09675_ team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\] net833 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[15\]
+ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout553_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ net914 _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08629__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net97 net2542 net891 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout720_A _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout818_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11703__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07508_ net991 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08488_ net919 _04273_ _04282_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__nor3_4
XANTENNA__09841__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12189__A0 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15949__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11004__A team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10450_ _05722_ net372 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] net713 _04790_ vssd1
+ vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12534__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _05094_ _05113_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nor2_1
XANTENNA__08801__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12120_ net284 net1962 net587 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12051_ net319 net2109 net530 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
Xhold380 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold391 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _04416_ _06304_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15329__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _04652_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_2
X_15810_ clknet_leaf_50_wb_clk_i _02261_ _00768_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout871 _04642_ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_8
X_16790_ net1344 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
Xfanout882 _04634_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15741_ clknet_leaf_114_wb_clk_i _02192_ _00699_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09144__A _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _06476_ net226 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16692__1246 vssd1 vssd1 vccd1 vccd1 _16692__1246/HI net1246 sky130_fd_sc_hd__conb_1
Xhold1080 net111 vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14985__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1091 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net249 net2311 net542 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XANTENNA__10675__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15672_ clknet_leaf_122_wb_clk_i _02123_ _00630_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12884_ team_02_WB.instance_to_wrap.top.pc\[7\] _05725_ vssd1 vssd1 vccd1 vccd1 _02918_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14623_ net1156 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
X_11835_ net594 _04578_ _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__or3_4
XFILLER_0_96_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11613__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ net1056 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
X_11766_ net360 net1963 net560 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09832__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10978__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ net1888 _03356_ _03357_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o21a_1
X_10717_ _06366_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nand2_1
X_14485_ net1120 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ net356 net2192 net571 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16224_ clknet_leaf_36_wb_clk_i _02669_ _01181_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13436_ net992 _03302_ _03316_ _03309_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09045__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10648_ _06251_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08399__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16155_ clknet_leaf_1_wb_clk_i net1472 _01113_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13367_ _03266_ _03268_ _03269_ _03210_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__or4b_1
XANTENNA__12444__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] net930 net591 vssd1
+ vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__a21o_1
X_15106_ clknet_leaf_47_wb_clk_i _01557_ _00064_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12318_ net269 net1725 net500 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__mux2_1
X_16086_ clknet_leaf_78_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[4\] _01044_
+ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__dfrtp_1
X_13298_ _03196_ _03205_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ net1156 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__inv_2
X_12249_ net316 net2600 net509 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09899__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ net341 _03679_ team_02_WB.instance_to_wrap.top.a1.dataIn\[13\] _03649_ vssd1
+ vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15939_ clknet_leaf_45_wb_clk_i _02390_ _00897_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10666__B1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _05124_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nor2_8
XANTENNA__08893__A team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10130__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ net991 _03418_ _04276_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__or3b_1
XANTENNA__08005__A1_N _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09391_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[22\] net867 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[22\]
+ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08342_ _04207_ _04215_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09823__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10969__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ _04146_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09036__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12354__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09229__A _04908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout670_A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16500__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07988_ _03841_ _03842_ _03860_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15621__CLK clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[14\] net879 net838 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12102__B _04428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _05320_ _05322_ _05324_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__or4_2
XFILLER_0_74_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10121__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] team_02_WB.instance_to_wrap.top.a1.instruction\[30\]
+ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__or4_1
X_09589_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[17\] net856 net795 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a22o_1
XANTENNA__12529__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11620_ net299 net2449 net577 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11551_ net423 _06794_ _07140_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ _05977_ _05978_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13359__C1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09027__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ net1022 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11482_ _06918_ _07082_ net393 vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__mux2_1
XANTENNA__08742__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ team_02_WB.START_ADDR_VAL_REG\[29\] _04356_ vssd1 vssd1 vccd1 vccd1 net213
+ sky130_fd_sc_hd__and2_1
XFILLER_0_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10433_ _06077_ _06085_ net399 _06072_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12264__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10188__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11385__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _03144_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10364_ _05656_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ net239 net2718 net586 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13083_ _07012_ net227 _03091_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__o211a_1
X_10295_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[1\] net777 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[1\]
+ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12034_ net359 net2030 net468 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XANTENNA__11399__A2_N _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11608__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16410__D team_02_WB.instance_to_wrap.top.ru.dmmload_co\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout690 _04468_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_8
X_16773_ net1327 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
X_13985_ net1143 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12936_ _02883_ _02884_ _02968_ _02881_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a31o_1
X_15724_ clknet_leaf_52_wb_clk_i _02175_ _00682_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ team_02_WB.instance_to_wrap.top.pc\[18\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _02901_ sky130_fd_sc_hd__and2_1
X_15655_ clknet_leaf_15_wb_clk_i _02106_ _00613_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12439__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14606_ net1194 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11818_ net269 net2569 net552 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09266__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15586_ clknet_leaf_49_wb_clk_i _02037_ _00544_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12798_ _07408_ _07419_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ net1025 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
X_11749_ net315 net1708 net562 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ net1143 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12682__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16207_ clknet_leaf_38_wb_clk_i _02652_ _01164_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[7\]
+ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[6\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or4b_1
XANTENNA__12174__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14399_ net1118 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16138_ clknet_leaf_129_wb_clk_i net1478 _01096_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13117__A2 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08960_ _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__inv_2
X_16069_ clknet_leaf_127_wb_clk_i _02520_ _01027_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15644__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _03748_ _03773_ _03750_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a21o_1
X_08891_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04429_ vssd1 vssd1
+ vccd1 vccd1 _04576_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07842_ _03717_ _03718_ _03716_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07773_ _03630_ _03635_ net350 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09512_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\] net815 net760 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[19\]
+ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10103__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[20\] net672 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[20\]
+ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a221o_1
XANTENNA__12349__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout349_A _07094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09257__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09374_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\] net660 net656 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\]
+ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _04194_ _04196_ _04187_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1160_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_A _07213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09009__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ _04127_ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15174__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12084__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08187_ _04030_ net224 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16691__1245 vssd1 vssd1 vccd1 vccd1 _16691__1245/HI net1245 sky130_fd_sc_hd__conb_1
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13108__A2 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10080_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[6\] net807 _05737_ _05739_
+ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13770_ net1013 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XANTENNA__09496__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _04993_ _06201_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12721_ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 _07348_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ clknet_leaf_36_wb_clk_i _01891_ _00398_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _07275_ _07276_ _07277_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__nor4_1
XANTENNA__09248__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11603_ net248 net2692 net578 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15517__CLK clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ clknet_leaf_20_wb_clk_i _01822_ _00329_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12583_ net283 net2621 net472 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
X_14322_ net1084 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11534_ net434 _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ net1131 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11465_ _05749_ net454 _06135_ _05748_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13204_ team_02_WB.START_ADDR_VAL_REG\[12\] net996 net932 vssd1 vssd1 vccd1 vccd1
+ net195 sky130_fd_sc_hd__a21o_1
X_10416_ _05134_ net372 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14184_ net1090 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ net416 _06605_ _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__a21o_1
XANTENNA__09420__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ net989 team_02_WB.instance_to_wrap.wb.curr_state\[0\] _04551_ _03404_ team_02_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10347_ _05978_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__and2_1
XANTENNA__14503__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13066_ _02913_ _02944_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10278_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12017_ net316 net2655 net470 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XANTENNA__10333__A2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ net152 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09487__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16756_ net1310 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
X_13968_ net1003 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15707_ clknet_leaf_118_wb_clk_i _02158_ _00665_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11581__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12169__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _02903_ _02952_ _02905_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a21oi_1
X_16687_ net1241 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13899_ net1030 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
XANTENNA__10478__A _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09239__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15638_ clknet_leaf_110_wb_clk_i _02089_ _00596_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15569_ clknet_leaf_17_wb_clk_i _02020_ _00527_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16442__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _03955_ _03984_ _03954_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09090_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\] net813 net854 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[29\]
+ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold72_A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08041_ _03886_ _03913_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold902 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 net108 vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[18\] vssd1 vssd1 vccd1
+ vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11214__A2_N net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold957 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _05646_ _05650_ _05652_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nor4_1
Xhold979 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08943_ team_02_WB.instance_to_wrap.top.a1.instruction\[23\] net930 _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\]
+ net740 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a221o_1
XANTENNA__08411__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08874_ _04273_ _04309_ _04320_ net940 team_02_WB.instance_to_wrap.top.a1.dataIn\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1006_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _03710_ _03715_ _03709_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout466_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07756_ _03408_ net350 _03608_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08557__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ _03562_ _03569_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_1656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12079__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09426_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[21\] net857 net833 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09357_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11711__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08308_ team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] _04165_ vssd1 vssd1 vccd1
+ vccd1 _04186_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\] net710 net641 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[24\]
+ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09650__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ _04071_ _04120_ _04097_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11250_ _06062_ _06087_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09402__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10201_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[3\] net881 net760 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\]
+ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ net317 net2658 net583 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XANTENNA__12542__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10132_ net595 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[5\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_101_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10063_ team_02_WB.instance_to_wrap.top.a1.instruction\[18\] net615 _04427_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__a22o_1
X_14940_ net999 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XANTENNA__11512__A1 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10315__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input27_A wbm_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ net1191 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16610_ clknet_leaf_67_wb_clk_i _02844_ _01483_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13822_ net1021 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13753_ net1062 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
X_16541_ clknet_leaf_129_wb_clk_i net1443 _01414_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10965_ _06605_ net413 net436 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and3b_1
XANTENNA__14993__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ team_02_WB.instance_to_wrap.top.pc\[1\] _04510_ vssd1 vssd1 vccd1 vccd1 _07332_
+ sky130_fd_sc_hd__nand2_1
X_13684_ net1039 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
X_16472_ clknet_leaf_99_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[7\] _01346_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10896_ net415 net436 _06540_ _06142_ net452 vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a32o_1
X_12635_ net410 _06531_ _07258_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__a211o_1
X_15423_ clknet_leaf_10_wb_clk_i _01874_ _00381_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11621__S net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15354_ clknet_leaf_120_wb_clk_i _01805_ _00312_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ net237 net2332 net474 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] net887 net907 team_02_WB.instance_to_wrap.top.pc\[4\]
+ _07114_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__a221o_1
X_14305_ net1144 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ clknet_leaf_115_wb_clk_i _01736_ _00243_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12497_ net360 net2056 net480 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__mux2_1
Xhold209 team_02_WB.instance_to_wrap.top.pc\[29\] vssd1 vssd1 vccd1 vccd1 net1607
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14236_ net1102 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _06330_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ net1108 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ net434 _06986_ _06989_ _06985_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__o211a_1
XANTENNA__10761__A _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _02930_ _03122_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__nor2_1
X_14098_ net1081 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10480__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _02948_ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07610_ _03499_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__or2_1
X_16808_ net1362 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
X_08590_ net976 _04376_ _04377_ _04382_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a311o_1
XFILLER_0_89_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire601_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ team_02_WB.instance_to_wrap.top.a1.dataIn\[25\] team_02_WB.instance_to_wrap.top.a1.dataIn\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__and2_1
XANTENNA__11267__B1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16739_ net1293 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
X_16690__1244 vssd1 vssd1 vccd1 vccd1 _16690__1244/HI net1244 sky130_fd_sc_hd__conb_1
XFILLER_0_53_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07472_ net996 vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15832__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09211_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[26\] net812 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[26\]
+ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09142_ net898 net613 _04630_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09632__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\] net706 net665 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15982__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08024_ _03893_ _03882_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__and2b_1
Xhold710 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\] vssd1 vssd1 vccd1
+ vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold743 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10671__A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold754 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15212__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16338__CLK clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11486__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[8\] net775 net842 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout583_A _04580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] net625 _04610_ vssd1
+ vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a21o_1
XANTENNA__13982__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08857_ net18 net950 _04555_ net1673 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout848_A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07808_ _03696_ _03698_ _03666_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21ai_1
X_08788_ _04551_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net925 vssd1 vssd1
+ vccd1 vccd1 _04552_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_93_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07739_ _03626_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__nor2_1
XANTENNA__13206__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ _05883_ net369 _06400_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09871__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09409_ _05077_ _05079_ _05081_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12537__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ team_02_WB.instance_to_wrap.top.pc\[11\] _06332_ vssd1 vssd1 vccd1 vccd1
+ _06333_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ net301 net1706 net490 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09623__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12351_ net268 net1933 net496 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_67_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11302_ net400 _06918_ _06915_ net409 vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ clknet_leaf_85_wb_clk_i _01521_ _00033_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_12282_ net316 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[18\] net506 vssd1
+ vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
XANTENNA__08750__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12780__B _05593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ net1076 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
X_11233_ net440 _06842_ _06855_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[16\]
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_120_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12272__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11164_ _06679_ _06790_ net383 vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14988__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[5\] net880 net876 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a22o_1
X_15972_ clknet_leaf_55_wb_clk_i _02423_ _00930_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11095_ _06722_ _06723_ _06726_ team_02_WB.instance_to_wrap.top.aluOut\[21\] net459
+ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__o32a_4
XFILLER_0_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ net1041 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
X_10046_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[6\] net730 net626 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 team_02_WB.instance_to_wrap.top.pc\[7\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[1\] vssd1 vssd1 vccd1 vccd1
+ net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[9\] vssd1 vssd1 vccd1
+ vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ net1166 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
X_13805_ net1134 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14785_ net1180 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
X_11997_ net2070 net343 net532 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ clknet_leaf_36_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[27\]
+ _01398_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13736_ net1096 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
X_10948_ _06143_ _06204_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16455_ clknet_leaf_81_wb_clk_i net1470 _01329_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12447__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ net1068 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
X_10879_ _06064_ _06093_ net387 vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15406_ clknet_leaf_42_wb_clk_i _01857_ _00364_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12618_ _06621_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__or2_1
X_16386_ clknet_leaf_73_wb_clk_i net1604 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13598_ net1020 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XANTENNA__09614__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15337_ clknet_leaf_24_wb_clk_i _01788_ _00295_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11421__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ net267 net2687 net464 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15235__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _04347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15268_ clknet_leaf_19_wb_clk_i _01719_ _00226_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12182__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14219_ net1030 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15199_ clknet_leaf_26_wb_clk_i _01650_ _00157_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09393__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout508 _07216_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_8
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout519 _07213_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_2
XANTENNA__14898__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] net797 net753 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[13\]
+ _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a221o_1
X_08711_ _04504_ net456 _04507_ net463 net741 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a221o_1
X_09691_ _05337_ _05355_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__nor2_1
XANTENNA__08353__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1095 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_4
X_08642_ net910 _04427_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__or2_4
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04366_ vssd1 vssd1 vccd1
+ vccd1 _04370_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07524_ team_02_WB.instance_to_wrap.top.a1.halfData\[2\] team_02_WB.instance_to_wrap.top.a1.halfData\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07455_ net976 vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16010__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12357__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13401__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[28\] net770 net834 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08959__A2 team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16160__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[30\] net818 net849 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[30\]
+ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ _03872_ net241 _03873_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout798_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15728__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12092__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold551 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold584 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09958_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[8\] net705 _05619_ vssd1
+ vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09136__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ net975 net976 _04406_ net974 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__and4b_1
X_09889_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[10\] net819 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ net293 net2279 net540 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
Xhold1273 team_02_WB.START_ADDR_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1284 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15108__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ net323 net2276 net548 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _06099_ _06104_ net365 vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14570_ net1036 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
X_11782_ net315 net2645 net558 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09844__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12775__B _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13521_ _03368_ _03369_ net885 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__and3b_1
X_10733_ _06382_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12267__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15258__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13452_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[11\] _03325_ vssd1 vssd1 vccd1
+ vccd1 _03326_ sky130_fd_sc_hd__and2_1
X_16240_ clknet_leaf_93_wb_clk_i _02678_ _01197_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input94_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ team_02_WB.instance_to_wrap.top.a1.instruction\[31\] net931 net591 vssd1
+ vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a21oi_1
X_12403_ net248 net2523 net491 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16171_ clknet_leaf_71_wb_clk_i _02617_ _01129_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ _03277_ _03283_ _03284_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10595_ team_02_WB.instance_to_wrap.top.pc\[22\] _06246_ vssd1 vssd1 vccd1 vccd1
+ _06247_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _07194_ _07214_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nand2b_1
X_15122_ clknet_leaf_15_wb_clk_i _01573_ _00080_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15053_ clknet_leaf_89_wb_clk_i _01504_ _00016_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_12265_ net353 net2385 net508 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07525__A_N team_02_WB.instance_to_wrap.top.a1.halfData\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10509__A2 _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ net1039 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
X_11216_ net909 _06838_ _06837_ net444 vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__a211o_1
X_12196_ net342 net1810 net516 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XANTENNA__10914__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ team_02_WB.instance_to_wrap.top.pc\[18\] _06337_ team_02_WB.instance_to_wrap.top.pc\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09127__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ net388 _06709_ _06710_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__o21ai_1
X_15955_ clknet_leaf_124_wb_clk_i _02406_ _00913_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14906_ net1164 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
X_10029_ _05683_ _05685_ _05687_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__or4_1
X_15886_ clknet_leaf_43_wb_clk_i _02337_ _00844_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10142__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14837_ net1193 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09835__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14768_ net1181 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16507_ clknet_leaf_129_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[10\]
+ _01381_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13719_ net1119 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XANTENNA__12177__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14699_ net1159 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16438_ clknet_leaf_99_wb_clk_i net1485 _01312_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16369_ clknet_leaf_74_wb_clk_i _02802_ _01261_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07795__A team_02_WB.instance_to_wrap.top.a1.dataIn\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _06780_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
Xfanout316 net318 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10905__C1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout327 net329 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlymetal6s2s_1
X_09812_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[12\] net815 net811 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[12\]
+ _05467_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a221o_1
Xfanout338 net340 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout349 _07094_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16785__1339 vssd1 vssd1 vccd1 vccd1 _16785__1339/HI net1339 sky130_fd_sc_hd__conb_1
XANTENNA__09118__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[13\] net736 net732 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[13\]
+ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout281_A _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[15\] net761 net757 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a22o_1
XANTENNA__08877__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08625_ net826 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net98 net1661 net894 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16526__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07507_ net4 net3 net2 net1 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__nor4_1
XFILLER_0_33_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12087__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _04320_ _04321_ _04324_ net751 net1687 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout713_A _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15550__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\] net737 net649 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10380_ _05156_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09039_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ net315 net1757 net529 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold370 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ net441 _06620_ _06639_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[24\]
+ sky130_fd_sc_hd__a21o_2
XANTENNA__12550__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout850 _04662_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09109__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout861 _04647_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout872 _04642_ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_2
Xfanout883 _04633_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_2
XANTENNA__16056__CLK clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout894 _04357_ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
X_15740_ clknet_leaf_48_wb_clk_i _02191_ _00698_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12952_ _02878_ _02971_ net229 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10124__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08868__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1070 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1081 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10675__A1 team_02_WB.instance_to_wrap.top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ net245 net2393 net542 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
Xhold1092 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
X_15671_ clknet_leaf_116_wb_clk_i _02122_ _00629_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12883_ _02915_ _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08983__B _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14622_ net1164 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11834_ team_02_WB.instance_to_wrap.top.a1.instruction\[10\] _04428_ team_02_WB.instance_to_wrap.top.a1.instruction\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__or3b_4
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11624__A0 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ net1061 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
XANTENNA__16408__D team_02_WB.instance_to_wrap.top.ru.dmmload_co\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ net352 net2024 net560 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13504_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\] _03356_ net873 vssd1
+ vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ _04804_ net368 vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14484_ net1050 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
X_11696_ net342 net2053 net568 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13377__B1 _03226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16223_ clknet_leaf_35_wb_clk_i _02668_ _01180_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\] _03301_ vssd1 vssd1 vccd1
+ vccd1 _03316_ sky130_fd_sc_hd__or2_1
X_10647_ _03402_ _06252_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ clknet_leaf_5_wb_clk_i _02600_ _01112_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
X_13366_ net987 _03212_ _03239_ team_02_WB.instance_to_wrap.top.a1.row1\[123\] vssd1
+ vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a22o_1
X_10578_ team_02_WB.instance_to_wrap.top.pc\[28\] _06228_ vssd1 vssd1 vccd1 vccd1
+ _06230_ sky130_fd_sc_hd__xnor2_1
X_15105_ clknet_leaf_130_wb_clk_i _01556_ _00063_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11552__A2_N net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ net323 net2273 net501 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
X_13297_ team_02_WB.instance_to_wrap.top.a1.halfData\[5\] _03174_ net995 vssd1 vssd1
+ vccd1 vccd1 _03205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16085_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[3\] _01043_
+ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09348__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15036_ net1149 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
X_12248_ net305 net2321 net511 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12179_ net288 net1848 net516 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XANTENNA__12460__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15938_ clknet_leaf_47_wb_clk_i _02389_ _00896_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10115__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16549__CLK clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15869_ clknet_leaf_114_wb_clk_i _02320_ _00827_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08893__B team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11804__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _00011_ _03419_ _04276_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[22\] net876 net839 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a22o_1
XANTENNA__09808__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08341_ _04209_ _04212_ _04216_ _04211_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15573__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ net2128 net937 net919 _04152_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11091__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14416__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09587__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08795__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__A_N team_02_WB.instance_to_wrap.top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09339__A2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12370__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout663_A _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09726_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[14\] net790 net774 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[14\]
+ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a221o_1
XANTENNA__10106__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[15\] net732 net636 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\]
+ _05325_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15916__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11714__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] team_02_WB.instance_to_wrap.top.a1.instruction\[28\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[27\] team_02_WB.instance_to_wrap.top.a1.instruction\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__or4_1
X_09588_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[17\] net780 net763 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13214__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08539_ net85 net1635 net893 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13071__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ _05934_ _06157_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__xor2_1
X_10501_ _05658_ _06150_ _06152_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__or4_1
XFILLER_0_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12545__S net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ _07002_ _07081_ net382 vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ team_02_WB.START_ADDR_VAL_REG\[28\] net61 net934 vssd1 vssd1 vccd1 vccd1
+ net212 sky130_fd_sc_hd__a21o_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09578__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ net384 _06084_ net393 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11385__A2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _03399_ _03137_ _03143_ net1184 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10363_ _05591_ _05613_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12102_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _04428_ _04578_ _04579_
+ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__or4_4
X_13082_ _07431_ _03092_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input57_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[1\] net853 net878 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12033_ net352 net2247 net468 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XANTENNA__12280__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14061__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A2 _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15446__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09750__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14996__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _04471_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout691 _04468_ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_2
X_16772_ net1326 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
X_13984_ net1071 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
X_15723_ clknet_leaf_22_wb_clk_i _02174_ _00681_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_12935_ _02884_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15596__CLK clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11624__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15654_ clknet_leaf_13_wb_clk_i _02105_ _00612_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12866_ team_02_WB.instance_to_wrap.top.pc\[18\] _06260_ vssd1 vssd1 vccd1 vccd1
+ _02900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ net1198 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11817_ net323 net2240 net552 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15585_ clknet_leaf_2_wb_clk_i _02036_ _00543_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12797_ _07407_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14536_ net1089 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ net304 net2440 net563 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16784__1338 vssd1 vssd1 vccd1 vccd1 _16784__1338/HI net1338 sky130_fd_sc_hd__conb_1
XFILLER_0_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12455__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ net1069 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ net287 net2189 net568 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16206_ clknet_leaf_7_wb_clk_i _02651_ _01163_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09569__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13418_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[5\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[4\]
+ _03301_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14398_ net1022 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08777__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16221__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16137_ clknet_leaf_1_wb_clk_i _02583_ _01095_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dfrtp_1
X_13349_ net2511 net895 _03253_ net992 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16068_ clknet_leaf_54_wb_clk_i _02519_ _01026_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08529__A0 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07910_ _03790_ _03791_ _03771_ _03779_ _03780_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a2111o_1
X_15019_ net1190 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12190__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ team_02_WB.instance_to_wrap.top.a1.row1\[101\] _03423_ vssd1 vssd1 vccd1
+ vccd1 _02532_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10336__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07841_ _03727_ _03728_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a21o_1
XANTENNA__09741__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15939__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07772_ _03635_ net350 vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__and2_1
X_09511_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[19\] net787 net776 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[20\] net720 net696 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09373_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[22\] net672 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08324_ _04199_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13119__A1_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08255_ net2461 net937 net919 _04136_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
XANTENNA__12365__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1153_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout509_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08186_ _04066_ _04068_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15469__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09980__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout878_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__S net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16511__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13209__B _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _05370_ _05372_ _05374_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__or4_4
X_10981_ _06042_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13292__A2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ team_02_WB.instance_to_wrap.top.a1.instruction\[19\] team_02_WB.instance_to_wrap.top.a1.instruction\[18\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[17\] team_02_WB.instance_to_wrap.top.a1.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12651_ _04700_ _05483_ _05522_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ net244 net2337 net578 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15370_ clknet_leaf_46_wb_clk_i _01821_ _00328_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09799__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ net269 net2289 net472 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12783__B _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ net1028 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XANTENNA__12275__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ net419 _06764_ _07124_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__inv_2
X_14252_ net1018 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ team_02_WB.START_ADDR_VAL_REG\[11\] net997 net933 vssd1 vssd1 vccd1 vccd1
+ net194 sky130_fd_sc_hd__a21o_1
X_10415_ _05094_ net367 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14183_ net1153 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_11395_ net399 _07003_ _07000_ net408 vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13134_ net6 _04341_ _04339_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__a21o_1
XANTENNA__10030__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _04502_ net370 vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__or2_1
XANTENNA__11619__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ team_02_WB.instance_to_wrap.top.pc\[12\] net945 _03079_ vssd1 vssd1 vccd1
+ vccd1 _01510_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10277_ net391 _05929_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__nor2_1
XANTENNA__10318__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ net304 net1916 net471 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XANTENNA__09723__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08931__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16824_ net152 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16755_ net1309 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ net1125 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XANTENNA__13283__A2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15706_ clknet_leaf_116_wb_clk_i _02157_ _00664_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10097__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ team_02_WB.instance_to_wrap.top.pc\[15\] _06268_ _02951_ vssd1 vssd1 vccd1
+ vccd1 _02952_ sky130_fd_sc_hd__a21oi_1
X_16686_ net1240 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__11294__B2 _06887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13898_ net1050 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15637_ clknet_leaf_115_wb_clk_i _02088_ _00595_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12849_ _02881_ _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ clknet_leaf_39_wb_clk_i _02019_ _00526_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08998__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ net1108 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12185__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ clknet_leaf_19_wb_clk_i _01950_ _00457_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08040_ _03892_ _03927_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap600 _05743_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold903 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold914 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold925 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10021__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold947 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09962__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold958 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\] net779 net759 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ _05638_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08942_ net977 net979 _04370_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a21o_1
XANTENNA__10309__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09714__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ net1559 _04564_ net825 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XANTENNA__08922__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ _03713_ _03711_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16117__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07755_ _03408_ _03608_ net350 vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout361_A _07170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07489__A0 team_02_WB.instance_to_wrap.top.a1.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__A0 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _03574_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[21\] net781 net761 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[21\]
+ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a221o_1
XANTENNA__13058__A1_N _07366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout626_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07978__A team_02_WB.instance_to_wrap.top.a1.dataIn\[8\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ _05012_ _05030_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__inv_2
X_09287_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] net653 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
XANTENNA__12095__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _04089_ _04090_ team_02_WB.instance_to_wrap.top.a1.dataIn\[4\] vssd1 vssd1
+ vccd1 vccd1 _04120_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10260__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _03944_ _04031_ _04051_ _04016_ _04029_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_82_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14604__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[3\] net784 net768 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10012__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ net444 _06783_ _06785_ team_02_WB.instance_to_wrap.top.aluOut\[18\] net460
+ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o32a_4
XFILLER_0_82_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09953__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _05782_ _05786_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__nor4_2
XFILLER_0_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09166__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10062_ _05712_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__nor2_4
XANTENNA__09705__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16783__1337 vssd1 vssd1 vccd1 vccd1 _16783__1337/HI net1337 sky130_fd_sc_hd__conb_1
X_14870_ net1186 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
XANTENNA__08748__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12778__B _05591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ net1105 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ clknet_leaf_128_wb_clk_i net1462 _01413_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10079__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13752_ net1056 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10964_ net401 _06604_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12703_ team_02_WB.instance_to_wrap.top.pc\[1\] _04510_ vssd1 vssd1 vccd1 vccd1 _07331_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16471_ clknet_leaf_99_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[6\] _01345_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[6\] sky130_fd_sc_hd__dfrtp_1
X_13683_ net1127 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
X_10895_ net400 _06539_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11902__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15422_ clknet_leaf_5_wb_clk_i _01873_ _00380_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _06880_ _07142_ _07260_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12776__A1 _05493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15353_ clknet_leaf_107_wb_clk_i _01804_ _00311_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12565_ team_02_WB.instance_to_wrap.top.a1.instruction\[11\] _07190_ _07205_ vssd1
+ vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__or3_4
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ net1070 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11516_ net914 _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__nor2_1
X_15284_ clknet_leaf_50_wb_clk_i _01735_ _00242_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _07153_ net2688 net480 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14235_ net1058 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
X_11447_ team_02_WB.instance_to_wrap.top.pc\[6\] _06329_ team_02_WB.instance_to_wrap.top.pc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10003__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__A1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ net1105 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XANTENNA__09944__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ net438 _06987_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08512__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10329_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[0\] net867 net847 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a22o_1
X_13117_ team_02_WB.instance_to_wrap.top.pc\[1\] _04510_ _02929_ vssd1 vssd1 vccd1
+ vccd1 _03122_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ net1078 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09157__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ team_02_WB.instance_to_wrap.top.pc\[14\] _06271_ vssd1 vssd1 vccd1 vccd1
+ _03065_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16807_ net1361 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
XANTENNA__15164__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14999_ net1186 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
X_07540_ team_02_WB.instance_to_wrap.top.a1.dataIn\[19\] team_02_WB.instance_to_wrap.top.a1.dataIn\[18\]
+ team_02_WB.instance_to_wrap.top.a1.dataIn\[17\] team_02_WB.instance_to_wrap.top.a1.dataIn\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11267__A1 team_02_WB.instance_to_wrap.top.a1.dataIn\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16738_ net1292 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XFILLER_0_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08407__A_N team_02_WB.instance_to_wrap.top.a1.halfData\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07471_ team_02_WB.instance_to_wrap.top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _03411_
+ sky130_fd_sc_hd__inv_2
X_16669_ net1224 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11812__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09210_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[26\] net866 net843 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ net614 vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.read_data2\[28\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09072_ team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[29\] net649 net633 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[29\]
+ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08023_ _03875_ _03877_ net241 vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__or3_1
Xhold700 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold711 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold722 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13192__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold733 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09935__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold744 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold766 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[4\] vssd1 vssd1 vccd1
+ vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09974_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1116_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08925_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[31\] net684 net676 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15507__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ net29 net950 net923 team_02_WB.instance_to_wrap.ramload\[2\] vssd1 vssd1
+ vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09253__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _03664_ _03697_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__or2_1
X_08787_ net984 team_02_WB.instance_to_wrap.top.ru.dmmWen vssd1 vssd1 vccd1 vccd1
+ _04551_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07738_ _03597_ _03625_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__and2_1
XANTENNA__09320__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ _03548_ _03553_ _03559_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11722__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[21\] net701 net652 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[21\]
+ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a221o_1
X_10680_ team_02_WB.instance_to_wrap.top.pc\[10\] team_02_WB.instance_to_wrap.top.pc\[9\]
+ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09339_ team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\] net812 net844 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[23\]
+ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12350_ net324 net2000 net496 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__D_N team_02_WB.instance_to_wrap.top.a1.instruction\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11301_ _06816_ _06917_ net382 vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12281_ net304 net2168 net507 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XANTENNA__12553__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14020_ net1141 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
X_11232_ net426 _06843_ _06846_ _06057_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__o221a_1
XANTENNA__09387__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09926__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11163_ _06735_ _06789_ net377 vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09139__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[5\] net855 net803 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ clknet_leaf_45_wb_clk_i _02422_ _00929_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11094_ net908 _06724_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14922_ net1001 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
X_10045_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[6\] net646 net618 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[6\]
+ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold60 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[7\] vssd1 vssd1 vccd1 vccd1
+ net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_02_WB.instance_to_wrap.top.pc\[16\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_02_WB.instance_to_wrap.top.pc\[8\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14853_ net1162 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
Xhold93 _02588_ vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ net1004 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14784_ net1177 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
X_11996_ net1749 net348 net534 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XANTENNA__09311__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16523_ clknet_leaf_35_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[26\]
+ _01397_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12997__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ net1153 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XANTENNA__12997__B2 _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10947_ _06143_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16454_ clknet_leaf_85_wb_clk_i net1589 _01328_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13666_ net1091 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10878_ _06142_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__xnor2_1
X_15405_ clknet_leaf_23_wb_clk_i _01856_ _00363_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12617_ _06703_ _06788_ _06957_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__or4_1
X_16385_ clknet_leaf_73_wb_clk_i _02816_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ net1080 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XANTENNA__10224__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15336_ clknet_leaf_57_wb_clk_i _01787_ _00294_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12548_ net324 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[16\] net464 vssd1
+ vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__mux2_1
XANTENNA__09090__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15267_ clknet_leaf_45_wb_clk_i _01718_ _00225_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12463__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net305 net2044 net482 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09378__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ net1037 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XANTENNA__09917__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15198_ clknet_leaf_12_wb_clk_i _01649_ _00156_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ net1073 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout509 _07216_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08710_ net975 net615 _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a21o_1
XANTENNA__11807__S net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11488__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1080 net1086 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_4
XANTENNA__09550__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08641_ team_02_WB.instance_to_wrap.top.i_ready net890 vssd1 vssd1 vccd1 vccd1 _04438_
+ sky130_fd_sc_hd__nand2_1
Xfanout1091 net1094 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12437__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04366_ vssd1 vssd1 vccd1
+ vccd1 _04369_ sky130_fd_sc_hd__nor2_1
XANTENNA__09302__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _03415_ _03416_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10999__B1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13323__A _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08417__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09124_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[28\] net813 net802 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a22o_1
XANTENNA__10215__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16782__1336 vssd1 vssd1 vccd1 vccd1 _16782__1336/HI net1336 sky130_fd_sc_hd__conb_1
XFILLER_0_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12881__B _05681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09055_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[30\] net863 net874 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a22o_1
XANTENNA__12373__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09369__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ _03874_ net241 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nor2_1
Xhold530 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold541 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold552 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold574 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold596 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[8\] net726 net718 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout860_A _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A _04340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__S net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08908_ _04388_ _04422_ _04433_ net581 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__and4_1
X_09888_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\] net771 net755 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\]
+ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__a221o_1
Xhold1230 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1241 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_02_WB.instance_to_wrap.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net2650
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ net17 net949 net923 team_02_WB.instance_to_wrap.ramload\[19\] vssd1 vssd1
+ vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
Xhold1263 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[9\] vssd1 vssd1 vccd1
+ vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1296 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ net322 net2026 net551 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _06092_ _06096_ net364 vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__mux2_1
XANTENNA__09711__A _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net303 net2477 net559 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11452__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13520_ team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[3\] _03366_
+ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10732_ _05378_ net369 vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13451_ net1175 _03324_ _03325_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__nor3_1
XFILLER_0_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ team_02_WB.instance_to_wrap.top.pc\[30\] _06223_ _06314_ vssd1 vssd1 vccd1
+ vccd1 _06315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12402_ net242 net2557 net489 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
X_16170_ clknet_leaf_71_wb_clk_i _02616_ _01128_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10206__A2 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11403__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_A wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10594_ net928 _05546_ net590 vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__a21o_2
XANTENNA__11403__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ net112 net896 net993 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09072__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15121_ clknet_leaf_17_wb_clk_i _01572_ _00079_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12333_ net233 net1887 net502 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__mux2_1
XANTENNA__12283__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14064__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15052_ clknet_leaf_99_wb_clk_i _01503_ _00015_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_12264_ net355 net2443 net511 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14003_ net1148 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
X_11215_ _06284_ _06286_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12195_ net348 net1715 net518 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__mux2_1
XANTENNA__10914__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15822__CLK clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _06258_ _06293_ _06294_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11627__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11077_ net384 _06599_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__or2_1
X_15954_ clknet_leaf_20_wb_clk_i _02405_ _00912_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09532__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ net1188 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
X_10028_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[7\] net821 net781 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[7\]
+ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a221o_1
X_15885_ clknet_leaf_32_wb_clk_i _02336_ _00843_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15972__CLK clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14836_ net1195 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12458__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ net1181 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11979_ net2055 net281 net534 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16729__1283 vssd1 vssd1 vccd1 vccd1 _16729__1283/HI net1283 sky130_fd_sc_hd__conb_1
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16506_ clknet_leaf_129_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[9\]
+ _01380_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15202__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13718_ net1084 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14698_ net1158 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ clknet_leaf_89_wb_clk_i net1493 _01311_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ net1078 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ clknet_leaf_74_wb_clk_i _02801_ _01260_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09063__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__A team_02_WB.instance_to_wrap.top.a1.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15352__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15319_ clknet_leaf_119_wb_clk_i _01770_ _00277_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12193__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16478__CLK clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16299_ clknet_leaf_98_wb_clk_i _02732_ _01242_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08810__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10905__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 _06780_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_1
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
X_09811_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[12\] net799 _05474_ _05476_
+ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a211o_1
XANTENNA__09771__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09742_ team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[13\] net692 net640 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10133__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\] net781 net777 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[15\]
+ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout274_A _06674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08624_ _04413_ _04417_ _04419_ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__nor4_1
XFILLER_0_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08555_ net99 net1579 net891 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12368__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11292__A1_N net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ team_02_WB.instance_to_wrap.top.pad.count\[1\] team_02_WB.instance_to_wrap.top.pad.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__and2_1
XFILLER_0_33_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08486_ _04317_ _04318_ net742 net751 net1572 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13988__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout706_A _04461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09054__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09107_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[28\] net729 net681 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\]
+ _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a221o_1
XANTENNA__16514__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08801__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09038_ _04712_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_8
XFILLER_0_60_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold360 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold371 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold382 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net428 _06621_ _06629_ net439 _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__a221o_1
Xhold393 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09762__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _04676_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
XANTENNA__13228__A net1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout851 _04662_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_8
Xfanout862 _04647_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_4
Xfanout873 _03337_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_2
Xfanout884 _03364_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_2
XANTENNA__09514__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout895 net896 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ team_02_WB.instance_to_wrap.top.pc\[30\] net943 net942 _02983_ vssd1 vssd1
+ vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1060 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11902_ net239 net2636 net542 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10675__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1082 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
X_15670_ clknet_leaf_109_wb_clk_i _02121_ _00628_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1093 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[25\] vssd1 vssd1 vccd1
+ vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08756__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12882_ team_02_WB.instance_to_wrap.top.pc\[8\] _05681_ vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14621_ net1167 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11833_ net235 net2098 net555 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
XANTENNA__12278__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14552_ net1054 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
X_11764_ net355 net2680 net563 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08057__A team_02_WB.instance_to_wrap.top.a1.dataIn\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13503_ _03356_ net873 _03355_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10715_ _04845_ net373 vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14483_ net1149 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11695_ net348 net2060 net569 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
XANTENNA__11910__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ clknet_leaf_38_wb_clk_i _02667_ _01179_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13434_ _03310_ _03315_ net1184 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a21oi_1
X_10646_ _06296_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09045__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ clknet_leaf_129_wb_clk_i net1504 _01111_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13365_ team_02_WB.instance_to_wrap.top.a1.row1\[3\] _03227_ _03230_ team_02_WB.instance_to_wrap.top.a1.row2\[43\]
+ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10577_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net930 net591 vssd1
+ vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a21o_1
XANTENNA__10060__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ clknet_leaf_9_wb_clk_i _01555_ _00062_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12316_ net321 net2212 net503 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16084_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[2\] _01042_
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__dfrtp_1
X_13296_ team_02_WB.instance_to_wrap.top.a1.halfData\[3\] _03174_ _03203_ _03204_
+ net995 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ net1151 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__inv_2
XANTENNA__08005__B1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ net298 net2209 net508 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12178_ net281 net1778 net518 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
X_11129_ _06524_ _06528_ net403 vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ clknet_leaf_1_wb_clk_i _02388_ _00895_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16781__1335 vssd1 vssd1 vccd1 vccd1 _16781__1335/HI net1335 sky130_fd_sc_hd__conb_1
X_15868_ clknet_leaf_48_wb_clk_i _02319_ _00826_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16150__CLK clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14819_ net1203 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ clknet_leaf_120_wb_clk_i _02250_ _00757_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08340_ _04201_ _04209_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08271_ _04142_ _04145_ _04149_ _04150_ _04140_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__a41o_2
XFILLER_0_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11091__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11820__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09036__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10051__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08547__A1 team_02_WB.START_ADDR_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15248__CLK clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07986_ _03835_ _03840_ _03860_ _03861_ _03838_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[14\] net794 net770 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout656_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[15\] net728 net692 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a22o_1
XANTENNA__07480__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ team_02_WB.instance_to_wrap.top.a1.instruction\[25\] net972 team_02_WB.instance_to_wrap.top.a1.instruction\[23\]
+ team_02_WB.instance_to_wrap.top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 _04404_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12098__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[17\] net776 net832 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout823_A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08538_ net86 net1602 net893 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08469_ net961 _04320_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11730__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ _05572_ _06146_ _06147_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__or3_1
XANTENNA__10290__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09027__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ _07037_ _07080_ net377 vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13230__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ _06080_ _06083_ net363 vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16822__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11031__A team_02_WB.instance_to_wrap.top.pc\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09983__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ team_02_WB.instance_to_wrap.top.lcd.nextState\[3\] _03137_ vssd1 vssd1 vccd1
+ vccd1 _03143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10362_ _05701_ _06014_ _05658_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16023__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12101_ net233 net1897 net526 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12561__S net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ _07431_ _03092_ net889 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a21oi_1
X_10293_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[1\] net813 net809 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14342__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ net354 net2096 net471 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
X_16728__1282 vssd1 vssd1 vccd1 vccd1 _16728__1282/HI net1282 sky130_fd_sc_hd__conb_1
Xhold190 team_02_WB.instance_to_wrap.top.a1.row1\[122\] vssd1 vssd1 vccd1 vccd1 net1588
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10345__A1 _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10896__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout670 _04477_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_8
Xfanout681 _04471_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_4
X_16771_ net1325 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
Xfanout692 _04467_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_6
X_13983_ net1130 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_15722_ clknet_leaf_43_wb_clk_i _02173_ _00680_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11905__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ _02967_ _02885_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15653_ clknet_leaf_128_wb_clk_i _02104_ _00611_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12865_ team_02_WB.instance_to_wrap.top.pc\[19\] _06257_ vssd1 vssd1 vccd1 vccd1
+ _02899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14604_ net1174 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
X_11816_ net322 net1997 net554 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15584_ clknet_leaf_12_wb_clk_i _02035_ _00542_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09266__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12796_ _05771_ _05768_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ net1136 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11747_ net296 net2132 net560 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11640__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14466_ net1091 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XANTENNA__10820__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11678_ net280 net1902 net568 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16205_ clknet_leaf_30_wb_clk_i _02650_ _01162_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13417_ net2411 _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ _06272_ _06278_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397_ net1081 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08777__B2 _04545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_36_wb_clk_i net1517 _01094_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap826 _04421_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ _03247_ _03249_ _03251_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16067_ clknet_leaf_45_wb_clk_i _02518_ _01025_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12471__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13279_ team_02_WB.instance_to_wrap.top.pad.keyCode\[3\] team_02_WB.instance_to_wrap.top.pad.keyCode\[2\]
+ team_02_WB.instance_to_wrap.top.pad.keyCode\[0\] team_02_WB.instance_to_wrap.top.pad.keyCode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__or4b_1
XFILLER_0_23_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15018_ net1190 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07840_ _03687_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07771_ _03627_ _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15540__CLK clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__S net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[19\] net792 net780 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[19\]
+ _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09081__A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _05114_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__inv_2
XANTENNA__13038__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[22\] net704 net692 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[22\]
+ _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a221o_1
XANTENNA__15690__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09257__A2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ _04183_ _04198_ _04178_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11064__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ _04127_ _04130_ _04134_ _04116_ _04113_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_69_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09009__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16046__CLK clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13210__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1146_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10024__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09965__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07475__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09717__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07969_ _03858_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nand2_4
XANTENNA__13277__B1 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[14\] net725 net653 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[14\]
+ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__a221o_1
X_10980_ _04993_ _06041_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__nor2_1
XANTENNA__09496__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09639_ team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[16\] net793 net837 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12650_ _05317_ _05357_ _05401_ _05441_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input104_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11601_ net239 net2469 net578 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12556__S net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ net323 net1935 net472 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14320_ net1016 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ net440 _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08208__B1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ net1030 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ net409 _06683_ _07064_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13202_ team_02_WB.START_ADDR_VAL_REG\[10\] net998 net934 vssd1 vssd1 vccd1 vccd1
+ net193 sky130_fd_sc_hd__a21o_1
X_16780__1334 vssd1 vssd1 vccd1 vccd1 _16780__1334/HI net1334 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08759__B2 _04536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _06065_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__nand2_1
XANTENNA__09956__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15413__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ net1140 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
X_11394_ _06917_ _07002_ net382 vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__mux2_1
XANTENNA__09420__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13133_ net1677 _03129_ _03126_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.nextHex\[3\]
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12291__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ _04510_ net898 _05996_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09708__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ _03074_ _03078_ _07366_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a21oi_1
X_10276_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ net296 net2508 net468 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16823_ net152 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11635__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13966_ net1114 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
X_16754_ net1308 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09487__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ clknet_leaf_107_wb_clk_i _02156_ _00663_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12917_ _02906_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16685_ net1239 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
X_13897_ net1024 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12848_ team_02_WB.instance_to_wrap.top.pc\[27\] _06235_ vssd1 vssd1 vccd1 vccd1
+ _02882_ sky130_fd_sc_hd__nor2_1
X_15636_ clknet_leaf_53_wb_clk_i _02087_ _00594_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09239__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ clknet_leaf_34_wb_clk_i _02018_ _00525_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12779_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__inv_2
XANTENNA__14247__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ net1109 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15498_ clknet_leaf_44_wb_clk_i _01949_ _00456_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14449_ net1029 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15093__CLK clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09947__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold904 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13087__A2_N net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap612 _05071_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09411__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__A1 _04846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold915 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16119_ clknet_leaf_64_wb_clk_i _02565_ _01077_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold937 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[5\] vssd1 vssd1 vccd1
+ vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold959 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[8\] net822 net862 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\]
+ _05651_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08941_ net977 net979 _04370_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ net959 _04306_ _04317_ net939 team_02_WB.instance_to_wrap.top.a1.dataIn\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07823_ _03713_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ _03637_ _03643_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09478__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ _03491_ _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout354_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1096_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[21\] net821 net841 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12884__B _05725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16727__1281 vssd1 vssd1 vccd1 vccd1 _16727__1281/HI net1281 sky130_fd_sc_hd__conb_1
X_09355_ _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout521_A _07212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _04177_ _04182_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09286_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\] net721 net629 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[24\]
+ _04963_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a221o_1
XANTENNA__09650__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ net2716 net936 net920 _04119_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09938__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08168_ _04030_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09402__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A _04362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_108_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15586__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16522__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ _03951_ _03956_ net225 _03957_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10130_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[5\] net867 net783 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[5\]
+ _05774_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ _05714_ _05716_ _05718_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__or4_2
XFILLER_0_41_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13236__A team_02_WB.instance_to_wrap.ramload\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13820_ net1123 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09469__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ net1111 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ net388 _06461_ _06465_ _06600_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12702_ net741 _07326_ _07329_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__or3b_1
X_16470_ clknet_leaf_99_wb_clk_i team_02_WB.instance_to_wrap.top.aluOut\[5\] _01344_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmaddr_co\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13682_ net1083 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
XANTENNA__08764__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10894_ net384 _06122_ _06535_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15421_ clknet_leaf_113_wb_clk_i _01872_ _00379_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12633_ net410 _06756_ _07165_ _07182_ net437 vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12286__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10595__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10236__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15352_ clknet_leaf_123_wb_clk_i _01803_ _00310_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12776__A2 _05502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12564_ net233 net1737 net465 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09641__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14303_ net1112 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11515_ _06328_ _07112_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15283_ clknet_leaf_3_wb_clk_i _01734_ _00241_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12495_ net356 net2202 net482 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ net1039 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ net429 _07036_ _07050_ net442 _07048_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[7\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA__10539__A1 _05215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ net1122 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
X_11377_ _05570_ net432 net454 _05572_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13116_ _07337_ _07341_ _07412_ net890 vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__o31ai_1
X_10328_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[0\] net791 net842 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[0\]
+ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a221o_1
X_14096_ net1003 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13047_ _07394_ _07438_ _07393_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21oi_1
X_10259_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[2\] net736 net716 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16806_ net1360 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_0_59_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14998_ net1187 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
X_16737_ net1291 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
X_13949_ net1054 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15459__CLK clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07470_ team_02_WB.instance_to_wrap.top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 _03410_
+ sky130_fd_sc_hd__inv_2
X_16668_ net1223 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_9_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15619_ clknet_leaf_42_wb_clk_i _02070_ _00577_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12196__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16599_ clknet_leaf_83_wb_clk_i _02833_ _01472_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _04815_ _04818_ _04820_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__nor4_2
XANTENNA__10936__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09093__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09632__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09071_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[29\] net729 net694 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a22o_1
XANTENNA__08840__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08022_ _03875_ _03894_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold712 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold723 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold745 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[27\] vssd1 vssd1 vccd1
+ vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08422__B _04277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold778 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ team_02_WB.instance_to_wrap.top.a1.instruction\[29\] net749 _05634_ vssd1
+ vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__o21a_2
XFILLER_0_106_1674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold789 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08924_ team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[31\] net664 net620 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1011_A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__B _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08855_ net32 net950 _04555_ net2650 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12782__A_N _05722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A _07193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _03630_ _03663_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09253__B _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ team_02_WB.instance_to_wrap.wb.curr_state\[1\] net6 vssd1 vssd1 vccd1 vccd1
+ _04550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07737_ _03624_ _03627_ _03622_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_A _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07668_ _03531_ _03555_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09871__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[21\] net672 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16517__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ _03470_ _03471_ _03453_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout903_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10218__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[23\] net852 net780 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09084__B1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08831__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[25\] net813 net855 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__A1_N team_02_WB.instance_to_wrap.top.a1.dataIn\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ _06871_ _06916_ net376 vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ net297 net2536 net504 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11231_ _05316_ net431 _06852_ _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_31_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12391__A0 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _06353_ _06358_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__nand2_1
XANTENNA__10941__A1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ net899 _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ clknet_leaf_49_wb_clk_i _02421_ _00928_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11093_ _06250_ _06251_ _06299_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__o21bai_1
XANTENNA_input32_A wbm_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\] net690 net657 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a22o_1
X_14921_ net1009 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[20\] vssd1 vssd1 vccd1 vccd1
+ net1448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold61 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[29\] vssd1 vssd1 vccd1 vccd1
+ net1459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08362__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1164 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
Xhold83 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[27\] vssd1 vssd1 vccd1
+ vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold94 team_02_WB.instance_to_wrap.top.a1.dataInTemp\[9\] vssd1 vssd1 vccd1 vccd1
+ net1492 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ net1013 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
X_14783_ net1183 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
X_11995_ net2270 net339 net534 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
XANTENNA_output119_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11913__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16522_ clknet_leaf_37_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[25\]
+ _01396_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13734_ net1142 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10946_ _04991_ _06042_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09862__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13665_ net1144 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
X_16453_ clknet_leaf_84_wb_clk_i net1558 _01327_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877_ _04910_ _06046_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10209__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15404_ clknet_leaf_52_wb_clk_i _01855_ _00362_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12616_ _07243_ _06977_ _06809_ _06730_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_52_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09075__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16384_ clknet_leaf_73_wb_clk_i _02815_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ net1123 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09614__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15335_ clknet_leaf_14_wb_clk_i _01786_ _00293_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12547_ net319 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[17\] net467 vssd1
+ vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ clknet_leaf_48_wb_clk_i _01717_ _00224_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ net296 net2679 net480 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ net1024 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11429_ net459 team_02_WB.instance_to_wrap.top.aluOut\[8\] _07034_ _06887_ vssd1
+ vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15197_ clknet_leaf_112_wb_clk_i _01648_ _00155_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14148_ net1094 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14079_ net1130 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
X_16726__1280 vssd1 vssd1 vccd1 vccd1 _16726__1280/HI net1280 sky130_fd_sc_hd__conb_1
XFILLER_0_83_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1070 net1072 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_4
XANTENNA__08353__A2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10696__B1 team_02_WB.instance_to_wrap.top.aluOut\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08640_ net462 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__inv_2
Xfanout1081 net1086 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1092 net1094 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_4
XANTENNA__15281__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__A2 _05797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08571_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] _04367_ vssd1 vssd1 vccd1
+ vccd1 _04368_ sky130_fd_sc_hd__and2_2
XFILLER_0_77_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11823__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07522_ team_02_WB.instance_to_wrap.top.pad.count\[0\] net991 vssd1 vssd1 vccd1 vccd1
+ _03416_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09853__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09066__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09605__A2 team_02_WB.instance_to_wrap.top.DUT.read_data2\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\] net866 net782 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08813__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14435__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09054_ team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[30\] net838 _04736_ _04737_
+ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08005_ _03894_ _03425_ net937 net2560 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a2bb2o_1
Xhold520 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12373__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold531 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[20\] vssd1 vssd1 vccd1
+ vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold542 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold553 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12912__A2 _05548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold575 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[12\] vssd1 vssd1 vccd1
+ vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[23\] vssd1 vssd1 vccd1
+ vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout686_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[8\] net673 net646 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[8\]
+ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__a221o_1
XANTENNA__07483__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ _04422_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__nand2_1
X_09887_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[10\] net787 net766 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__a22o_1
XANTENNA__12676__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_02_WB.instance_to_wrap.top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 net2618
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ net19 net947 net921 net1664 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__o22a_1
Xhold1242 team_02_WB.instance_to_wrap.top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 net2640
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\] vssd1 vssd1 vccd1
+ vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1264 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1286 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[2\] vssd1 vssd1 vccd1
+ vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ net1605 net955 net926 _04541_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
Xhold1297 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15774__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10800_ net394 _06445_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11780_ net297 net2340 net556 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09844__A2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A team_02_WB.instance_to_wrap.top.a1.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13233__B net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ _05421_ net374 vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16825__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[10\] team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[9\]
+ _03321_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10662_ _06226_ _06313_ _06224_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ net237 net2632 net489 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11969__A team_02_WB.instance_to_wrap.top.a1.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08804__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _03279_ _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nor2_1
XANTENNA__12564__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ team_02_WB.instance_to_wrap.top.pc\[23\] _04629_ vssd1 vssd1 vccd1 vccd1
+ _06245_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15120_ clknet_leaf_36_wb_clk_i _01571_ _00078_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12332_ net359 net2378 net500 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XANTENNA__10592__B _04629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15051_ clknet_leaf_90_wb_clk_i _01502_ _00014_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12263_ net343 net2036 net510 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14002_ net1082 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
X_11214_ team_02_WB.instance_to_wrap.top.a1.dataIn\[16\] net458 _06836_ net914 vssd1
+ vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_107_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12194_ net337 net2649 net518 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
XANTENNA__10914__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__S net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11145_ net441 _06755_ _06773_ net429 _06771_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.aluOut\[19\]
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11076_ _06648_ _06708_ net376 vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__mux2_1
X_15953_ clknet_leaf_17_wb_clk_i _02404_ _00911_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11209__A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ net1191 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
X_10027_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[7\] net869 net814 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a22o_1
XANTENNA__10113__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15884_ clknet_leaf_23_wb_clk_i _02335_ _00842_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10142__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14835_ net1166 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11643__S net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09296__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14766_ net1183 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11978_ net2697 net271 net535 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XANTENNA__08518__A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ clknet_leaf_0_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[8\]
+ _01379_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13717_ net1119 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
X_10929_ net387 _06379_ net394 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__o21a_1
X_14697_ net1157 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ clknet_leaf_91_wb_clk_i net1705 _01310_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13648_ net1016 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10783__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12474__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16367_ clknet_leaf_102_wb_clk_i _02800_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13579_ net1170 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10602__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__B _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15318_ clknet_leaf_109_wb_clk_i _01769_ _00276_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16298_ clknet_leaf_98_wb_clk_i _02731_ _01241_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15249_ clknet_leaf_17_wb_clk_i _01700_ _00207_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout307 _06975_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
XANTENNA__10905__B2 team_02_WB.instance_to_wrap.top.a1.dataIn\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09810_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[12\] net859 net880 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[12\]
+ _05475_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a221o_1
XANTENNA__11818__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout318 _06806_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_103_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout329 _07015_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
X_09741_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[13\] net680 _05407_ vssd1
+ vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15797__CLK clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09672_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[15\] net817 net814 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__a22o_1
XANTENNA__10133__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07534__B1 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ _04371_ _04418_ _04414_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08554_ net100 net1663 net891 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XANTENNA__09287__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09826__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07505_ net1646 net2743 net969 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12830__A1 _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08485_ _04314_ _04315_ net742 net751 net1658 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12384__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14165__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16422__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07478__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[28\] net733 net653 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09037_ _04714_ _04716_ _04718_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold350 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09211__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[13\] vssd1 vssd1 vccd1
+ vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_02_WB.instance_to_wrap.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net1781
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout830 net832 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
Xfanout841 _04672_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_8
Xfanout852 _04662_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13228__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ team_02_WB.instance_to_wrap.top.DUT.register\[14\]\[9\] net787 net779 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[9\]
+ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__a221o_1
Xfanout863 _04647_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_8
Xfanout874 _04668_ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_8
Xfanout885 _03364_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__dlymetal6s2s_1
X_12950_ _02872_ _02981_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__o21ai_1
Xfanout896 _03141_ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_2
Xhold1050 team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10124__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1061 team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net594 _07190_ _07199_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or3_4
XFILLER_0_38_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1072 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ team_02_WB.instance_to_wrap.top.pc\[8\] _05681_ vssd1 vssd1 vccd1 vccd1 _02915_
+ sky130_fd_sc_hd__nand2_1
Xhold1094 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__C _05929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14620_ net1167 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
X_11832_ net358 net1823 net552 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09278__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ net1112 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11763_ net342 net2564 net560 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10714_ net406 _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\] team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[12\]
+ _03353_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__and3_1
XANTENNA__08772__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14482_ net1084 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
X_11694_ net338 net2222 net569 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16221_ clknet_leaf_38_wb_clk_i _02666_ _01178_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13433_ _03301_ _03314_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__or2_1
X_10645_ team_02_WB.instance_to_wrap.top.pc\[20\] _06252_ vssd1 vssd1 vccd1 vccd1
+ _06297_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12294__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16152_ clknet_leaf_27_wb_clk_i net1513 _01110_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13364_ team_02_WB.instance_to_wrap.top.a1.row2\[27\] _03237_ _03238_ team_02_WB.instance_to_wrap.top.a1.row2\[35\]
+ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__a22o_1
X_10576_ team_02_WB.instance_to_wrap.top.a1.instruction\[28\] net930 net591 vssd1
+ vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12315_ net316 net2535 net500 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__mux2_1
X_15103_ clknet_leaf_8_wb_clk_i _01554_ _00061_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16083_ clknet_leaf_79_wb_clk_i team_02_WB.instance_to_wrap.top.a1.nextHex\[1\] _01041_
+ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.hexop\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13295_ _03180_ _03189_ _03193_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__or3_1
XFILLER_0_107_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14803__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ net1154 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
X_12246_ net288 net2317 net508 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16645__1216 vssd1 vssd1 vccd1 vccd1 _16645__1216/HI net1216 sky130_fd_sc_hd__conb_1
XFILLER_0_23_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_91_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11638__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12177_ net274 net1831 net518 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11128_ _06756_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__inv_2
X_16635__1383 vssd1 vssd1 vccd1 vccd1 net1383 _16635__1383/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15936_ clknet_leaf_7_wb_clk_i _02387_ _00894_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11059_ _04416_ _06301_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nor2_1
XANTENNA__10115__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12469__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15867_ clknet_leaf_104_wb_clk_i _02318_ _00825_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14818_ net1203 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09808__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15798_ clknet_leaf_110_wb_clk_i _02249_ _00756_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14749_ net1182 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08270_ _04145_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nand3_1
XFILLER_0_80_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16419_ clknet_leaf_60_wb_clk_i team_02_WB.instance_to_wrap.top.ru.dmmload_co\[18\]
+ _01293_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.dataIn\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08795__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__B1 _06629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07985_ _03863_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749__1303 vssd1 vssd1 vccd1 vccd1 _16749__1303/HI net1303 sky130_fd_sc_hd__conb_1
X_09724_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[14\] net870 _05381_ _05391_
+ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11303__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10106__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__B _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09655_ team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[15\] net616 _05323_ vssd1
+ vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a21o_1
XANTENNA__12379__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout551_A _07200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10688__A team_02_WB.instance_to_wrap.top.pc\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ team_02_WB.instance_to_wrap.top.a1.instruction\[6\] team_02_WB.instance_to_wrap.top.a1.instruction\[3\]
+ _04358_ net979 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _05247_ _05256_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__nor2_4
XFILLER_0_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ net87 net1637 net892 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08468_ team_02_WB.instance_to_wrap.top.a1.dataInTemp\[0\] _04277_ vssd1 vssd1 vccd1
+ vccd1 _04321_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15812__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16705__1259 vssd1 vssd1 vccd1 vccd1 _16705__1259/HI net1259 sky130_fd_sc_hd__conb_1
X_08399_ net1709 net935 net918 _04267_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ _06081_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10361_ _05747_ _06013_ _05703_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15962__CLK clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ net359 net1839 net525 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ _07403_ _07404_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__nor2_1
X_10292_ _05941_ _05943_ _05944_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11458__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net345 net2376 net469 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold180 team_02_WB.instance_to_wrap.top.a1.data\[9\] vssd1 vssd1 vccd1 vccd1 net1578
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_02_WB.instance_to_wrap.top.pc\[21\] vssd1 vssd1 vccd1 vccd1 net1589
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10345__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A3 _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 _04480_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout671 _04477_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_4
X_16770_ net1324 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
Xfanout682 _04471_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_6
XANTENNA__09499__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13982_ net1021 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
Xfanout693 _04467_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
X_15721_ clknet_leaf_24_wb_clk_i _02172_ _00679_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12933_ team_02_WB.instance_to_wrap.top.pc\[25\] _06242_ _02966_ vssd1 vssd1 vccd1
+ vccd1 _02967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12289__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15652_ clknet_leaf_54_wb_clk_i _02103_ _00610_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12864_ team_02_WB.instance_to_wrap.top.pc\[20\] _06255_ vssd1 vssd1 vccd1 vccd1
+ _02898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14603_ net1178 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
X_11815_ net315 net2665 net553 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ _07409_ _07416_ _07418_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__o21a_1
X_15583_ clknet_leaf_8_wb_clk_i _02034_ _00541_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11921__S net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14534_ net1141 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11746_ net290 net2052 net560 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09671__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14465_ net1143 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
X_11677_ net273 net1832 net571 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ clknet_leaf_29_wb_clk_i _02649_ _01161_ vssd1 vssd1 vccd1 vccd1 team_02_WB.START_ADDR_VAL_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10628_ _06269_ _06279_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nand2_1
X_13416_ team_02_WB.instance_to_wrap.top.lcd.cnt_20ms\[3\] _03300_ vssd1 vssd1 vccd1
+ vccd1 _03301_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09423__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14396_ net1110 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16135_ clknet_leaf_129_wb_clk_i net1515 _01093_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11230__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ team_02_WB.instance_to_wrap.top.a1.row1\[17\] _03222_ _03223_ team_02_WB.instance_to_wrap.top.a1.row1\[9\]
+ _03142_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10559_ _04785_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09627__A _05296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16066_ clknet_leaf_47_wb_clk_i _02517_ _01024_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13278_ _03181_ _03184_ _03185_ _03188_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15017_ net1190 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__inv_2
XANTENNA__13149__A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net347 net2330 net514 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap614_A _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12988__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _03598_ _03626_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15919_ clknet_leaf_33_wb_clk_i _02370_ _00877_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12199__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _05094_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[22\] net685 net648 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08322_ _04178_ _04183_ _04198_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09662__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12739__A_N team_02_WB.instance_to_wrap.top.i_ready vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08253_ _04127_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15985__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ _04019_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15215__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08441__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10690__B team_02_WB.instance_to_wrap.top.pc\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A _04674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16610__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _03800_ _03825_ _03853_ _03799_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a22o_4
XANTENNA__10910__S net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09707_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[14\] net700 net638 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ _03772_ _03782_ _03788_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_134_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09638_ team_02_WB.instance_to_wrap.top.DUT.register\[30\]\[16\] net821 net841 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09569_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[17\] net683 net643 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[17\]
+ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11600_ net594 _04579_ _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16644__1215 vssd1 vssd1 vccd1 vccd1 _16644__1215/HI net1215 sky130_fd_sc_hd__conb_1
XANTENNA__11741__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ net320 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[17\] net475 vssd1
+ vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ _06007_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__or2_1
XANTENNA__13241__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14250_ net1051 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XANTENNA__08208__A1 team_02_WB.instance_to_wrap.top.a1.row2\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16634__1382 vssd1 vssd1 vccd1 vccd1 net1382 _16634__1382/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11462_ net418 _06682_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09405__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ team_02_WB.START_ADDR_VAL_REG\[9\] net997 net932 vssd1 vssd1 vccd1 vccd1
+ net223 sky130_fd_sc_hd__a21o_1
XANTENNA__08759__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _05052_ net372 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14181_ net1073 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XANTENNA__12572__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11393_ _06959_ _07001_ net376 vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__mux2_1
X_13132_ team_02_WB.instance_to_wrap.top.a1.hexop\[1\] team_02_WB.instance_to_wrap.top.a1.hexop\[2\]
+ team_02_WB.instance_to_wrap.top.a1.hexop\[3\] vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or3_1
XANTENNA_input62_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _04510_ net898 _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ net230 _03076_ _03077_ _07436_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__o2bb2a_1
X_10275_ net391 _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nand2_2
XANTENNA__10318__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net287 net1943 net468 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11916__S net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16822_ net152 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08931__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16753_ net1307 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ net1135 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15704_ clknet_leaf_126_wb_clk_i _02155_ _00662_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12916_ team_02_WB.instance_to_wrap.top.pc\[14\] _06271_ _02949_ vssd1 vssd1 vccd1
+ vccd1 _02950_ sky130_fd_sc_hd__a21o_1
X_16684_ net1238 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__09892__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ net1100 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
X_15635_ clknet_leaf_125_wb_clk_i _02086_ _00593_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12847_ team_02_WB.instance_to_wrap.top.pc\[27\] _06235_ vssd1 vssd1 vccd1 vccd1
+ _02881_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ clknet_leaf_40_wb_clk_i _02017_ _00524_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09644__B1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12778_ _05593_ _05591_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14517_ net1120 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08998__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ net346 net2083 net565 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
X_15497_ clknet_leaf_31_wb_clk_i _01948_ _00455_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16748__1302 vssd1 vssd1 vccd1 vccd1 _16748__1302/HI net1302 sky130_fd_sc_hd__conb_1
XFILLER_0_126_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14448_ net1006 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12482__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14379_ net1026 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
Xhold905 team_02_WB.instance_to_wrap.top.DUT.register\[21\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[14\] vssd1 vssd1 vccd1
+ vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ clknet_leaf_63_wb_clk_i _02564_ _01076_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.ramload\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold938 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[17\] vssd1 vssd1 vccd1
+ vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15388__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ net580 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__inv_2
X_16049_ clknet_leaf_18_wb_clk_i _02500_ _01007_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10309__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ net1555 _04563_ net825 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ _03653_ _03680_ _03704_ _03712_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__11826__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13607__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08922__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16704__1258 vssd1 vssd1 vccd1 vccd1 _16704__1258/HI net1258 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07753_ _03578_ _03639_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07684_ _03524_ _03530_ _03556_ _03526_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[21\] net845 net765 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[21\]
+ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14438__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1089_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ net900 team_02_WB.instance_to_wrap.top.DUT.read_data2\[23\] net592 vssd1
+ vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07978__C _03859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ _04182_ _04177_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09285_ team_02_WB.instance_to_wrap.top.DUT.register\[23\]\[24\] net733 net625 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout514_A _07215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ _04107_ _04115_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__a21o_2
XFILLER_0_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ _04050_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__nand2_1
XANTENNA__12392__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07486__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ _03955_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09166__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10060_ team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[6\] net705 net622 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[6\]
+ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11736__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11037__A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ net413 _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ net1106 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09874__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _07327_ _07328_ team_02_WB.instance_to_wrap.top.aluOut\[31\] vssd1 vssd1
+ vccd1 vccd1 _07329_ sky130_fd_sc_hd__mux2_1
XANTENNA__12567__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ net1070 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
X_10893_ _06132_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15420_ clknet_leaf_49_wb_clk_i _01871_ _00378_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12632_ _07105_ _07259_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__nand2_1
XANTENNA__08429__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15351_ clknet_leaf_119_wb_clk_i _01802_ _00309_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12563_ net360 net2348 net467 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14302_ net1023 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
X_11514_ team_02_WB.instance_to_wrap.top.pc\[3\] team_02_WB.instance_to_wrap.top.pc\[2\]
+ team_02_WB.instance_to_wrap.top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12494_ net343 net2377 net480 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
X_15282_ clknet_leaf_15_wb_clk_i _01733_ _00240_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08780__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13398__S _03137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14233_ net1059 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
X_11445_ _06014_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14164_ net1039 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ net422 _06576_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ team_02_WB.instance_to_wrap.top.pc\[3\] net945 net942 _03120_ vssd1 vssd1
+ vccd1 vccd1 _01501_ sky130_fd_sc_hd__a22o_1
X_10327_ team_02_WB.instance_to_wrap.top.DUT.register\[7\]\[0\] net871 net881 team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14095_ net1129 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ team_02_WB.instance_to_wrap.top.pc\[15\] net946 net942 _03063_ vssd1 vssd1
+ vccd1 vccd1 _01513_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15680__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[2\] net628 net616 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[2\]
+ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11646__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[3\] net848 net840 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__a22o_1
XANTENNA__10172__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16805_ net1359 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XANTENNA__16036__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ net1187 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16736_ net1290 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
X_13948_ net1097 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XANTENNA__09865__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11672__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16667_ net1222 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__12477__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ net1111 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13162__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15618_ clknet_leaf_49_wb_clk_i _02069_ _00576_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16186__CLK clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16598_ clknet_leaf_75_wb_clk_i _02832_ _01471_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15549_ clknet_leaf_111_wb_clk_i _02000_ _00507_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09070_ _04746_ _04748_ _04750_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__or4_4
XFILLER_0_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08840__B2 team_02_WB.instance_to_wrap.ramload\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ _03902_ _03907_ _03897_ _03899_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11410__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold724 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_02_WB.instance_to_wrap.top.DUT.register\[29\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold746 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[24\] vssd1 vssd1 vccd1
+ vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold757 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[19\] vssd1 vssd1 vccd1
+ vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold768 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold779 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net463 _04509_ _05545_ net456 net741 vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a221o_1
XANTENNA__09148__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16643__1214 vssd1 vssd1 vccd1 vccd1 _16643__1214/HI net1214 sky130_fd_sc_hd__conb_1
X_08923_ team_02_WB.instance_to_wrap.top.DUT.register\[12\]\[31\] net736 net668 team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _06753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net33 net948 net922 team_02_WB.instance_to_wrap.ramload\[4\] vssd1 vssd1
+ vccd1 vccd1 _02549_ sky130_fd_sc_hd__o22a_1
XANTENNA__10163__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07805_ _03678_ _03679_ _03670_ _03672_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a211o_1
X_08785_ net1655 net958 net926 _04549_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a22o_1
X_16633__1381 vssd1 vssd1 vccd1 vccd1 net1381 _16633__1381/LO sky130_fd_sc_hd__conb_1
XANTENNA_fanout464_A _07225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _03597_ _03599_ _03625_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08865__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12895__B _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _03524_ _03556_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__xor2_2
XANTENNA__12387__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout729_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[21\] net640 _05080_ vssd1
+ vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__a21o_1
X_07598_ _03483_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__and2_1
XANTENNA__09608__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15553__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09337_ team_02_WB.instance_to_wrap.top.DUT.register\[19\]\[23\] net868 net816 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09268_ team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[25\] net771 net760 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[25\]
+ _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08219_ _04069_ _04099_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09199_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[26\] net696 net624 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11230_ _05318_ net455 net446 _05317_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09387__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16819__1373 vssd1 vssd1 vccd1 vccd1 _16819__1373/HI net1373 sky130_fd_sc_hd__conb_1
X_11161_ _05238_ _06190_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ team_02_WB.instance_to_wrap.top.a1.instruction\[26\] _04424_ _05770_ vssd1
+ vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__o21a_2
XFILLER_0_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11092_ _06250_ _06251_ _06299_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10043_ _05701_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor2_2
X_14920_ net1007 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XANTENNA__10154__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[17\] vssd1 vssd1 vccd1 vccd1
+ net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[6\] vssd1 vssd1 vccd1 vccd1
+ net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[31\] vssd1 vssd1 vccd1 vccd1
+ net1460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input25_A wbm_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ net1158 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
Xhold73 team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmstore\[22\] vssd1 vssd1 vccd1
+ vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
X_16747__1301 vssd1 vssd1 vccd1 vccd1 _16747__1301/HI net1301 sky130_fd_sc_hd__conb_1
Xhold84 _02606_ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_02_WB.instance_to_wrap.top.pc\[4\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ net1050 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09847__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14782_ net1182 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
X_11994_ net1808 net334 net532 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XANTENNA__09311__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ clknet_leaf_7_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[24\]
+ _01395_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13733_ net1089 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
XANTENNA__12297__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ net260 net1849 net585 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16452_ clknet_leaf_82_wb_clk_i net1483 _01326_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13664_ net1075 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10876_ net252 net2481 net583 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ clknet_leaf_22_wb_clk_i _01854_ _00361_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _06997_ _07242_ _07016_ _06843_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__nand4b_1
XANTENNA__11406__B1 _06886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16383_ clknet_leaf_73_wb_clk_i _02814_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pad.button_control.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ net1033 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14806__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15334_ clknet_leaf_13_wb_clk_i _01785_ _00292_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08822__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ net316 net1756 net466 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16703__1257 vssd1 vssd1 vccd1 vccd1 _16703__1257/HI net1257 sky130_fd_sc_hd__conb_1
X_15265_ clknet_leaf_129_wb_clk_i _01716_ _00223_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12477_ net289 net2214 net480 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 _07286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14216_ net1096 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XANTENNA__09378__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ team_02_WB.instance_to_wrap.top.pc\[8\] net907 _06886_ team_02_WB.instance_to_wrap.top.a1.dataIn\[8\]
+ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__a221o_1
X_15196_ clknet_leaf_49_wb_clk_i _01647_ _00154_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ net1073 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11359_ team_02_WB.instance_to_wrap.top.pc\[11\] _06332_ vssd1 vssd1 vccd1 vccd1
+ _06971_ sky130_fd_sc_hd__nor2_1
XANTENNA__08050__A2 _03933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14078_ net1022 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ _02902_ _02953_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10145__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15426__CLK clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1066 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
XANTENNA__09550__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10696__B2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1086 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_4
Xfanout1093 net1094 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_4
X_08570_ net979 _04366_ net978 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_83_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07521_ net1751 _03415_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16719_ net1273 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__09302__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15576__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10999__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11405__A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _04794_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__nor2_8
XFILLER_0_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12070__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__A _04510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[30\] net858 net777 team_02_WB.instance_to_wrap.top.DUT.register\[20\]\[30\]
+ _04728_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08004_ _03882_ _03891_ _03893_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09369__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[21\] vssd1 vssd1 vccd1
+ vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold521 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[8\] vssd1 vssd1 vccd1
+ vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold532 team_02_WB.instance_to_wrap.top.DUT.register\[9\]\[22\] vssd1 vssd1 vccd1
+ vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[0\] vssd1 vssd1 vccd1
+ vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 team_02_WB.instance_to_wrap.top.DUT.register\[26\]\[1\] vssd1 vssd1 vccd1
+ vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold576 team_02_WB.instance_to_wrap.top.DUT.register\[13\]\[28\] vssd1 vssd1 vccd1
+ vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold587 team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[26\] vssd1 vssd1 vccd1
+ vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[10\] vssd1 vssd1 vccd1
+ vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ team_02_WB.instance_to_wrap.top.DUT.register\[31\]\[8\] net698 net666 team_02_WB.instance_to_wrap.top.DUT.register\[24\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a22o_1
X_08906_ _04430_ _04586_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nor3_1
XFILLER_0_77_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09886_ team_02_WB.instance_to_wrap.top.DUT.register\[16\]\[10\] net803 net831 team_02_WB.instance_to_wrap.top.DUT.register\[17\]\[10\]
+ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a221o_1
Xhold1210 team_02_WB.instance_to_wrap.top.DUT.register\[1\]\[30\] vssd1 vssd1 vccd1
+ vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1221 team_02_WB.instance_to_wrap.top.DUT.register\[4\]\[15\] vssd1 vssd1 vccd1
+ vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[31\] vssd1 vssd1 vccd1
+ vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1243 team_02_WB.instance_to_wrap.top.DUT.register\[18\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net20 net949 net923 net1689 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1254 team_02_WB.instance_to_wrap.top.DUT.register\[2\]\[29\] vssd1 vssd1 vccd1
+ vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A _04664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1265 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15919__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1276 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[11\] vssd1 vssd1 vccd1
+ vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[6\] vssd1 vssd1 vccd1
+ vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 team_02_WB.instance_to_wrap.top.DUT.register\[15\]\[3\] vssd1 vssd1 vccd1
+ vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11018__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ team_02_WB.instance_to_wrap.top.ru.m1.prev_dmmaddr\[8\] team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[8\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__mux2_2
X_07719_ team_02_WB.instance_to_wrap.top.a1.dataIn\[15\] _03541_ _03582_ vssd1 vssd1
+ vccd1 vccd1 _03610_ sky130_fd_sc_hd__or3_1
XANTENNA__13102__A1_N net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16528__D team_02_WB.instance_to_wrap.top.DUT.read_data2\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08699_ net747 _04449_ _04466_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08608__B team_02_WB.instance_to_wrap.top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ net384 _06372_ _06380_ net399 vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ _06312_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12400_ _04576_ _07188_ _07199_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ team_02_WB.instance_to_wrap.top.a1.row2\[12\] _03206_ _03280_ _03273_ team_02_WB.instance_to_wrap.top.a1.row1\[108\]
+ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__a32o_1
X_10592_ team_02_WB.instance_to_wrap.top.pc\[23\] _04629_ vssd1 vssd1 vccd1 vccd1
+ _06244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ net353 net2320 net501 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12262_ net349 net2069 net510 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
X_15050_ clknet_leaf_90_wb_clk_i _01501_ _00013_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.pc\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11213_ _06336_ _06835_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__or2_1
X_14001_ net1030 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XANTENNA__12580__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ net334 net2646 net516 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10914__A2 _06323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11144_ _06193_ _06772_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__and2_1
XANTENNA__09780__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15952_ clknet_leaf_39_wb_clk_i _02403_ _00910_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11075_ _06066_ _06068_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14903_ net1187 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
X_10026_ team_02_WB.instance_to_wrap.top.DUT.register\[11\]\[7\] net817 net761 team_02_WB.instance_to_wrap.top.DUT.register\[22\]\[7\]
+ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a221o_1
XANTENNA__09532__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15599__CLK clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ clknet_leaf_21_wb_clk_i _02334_ _00841_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10113__B _05771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__S net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14834_ net1161 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14765_ net1181 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11977_ net2448 net275 net533 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
X_16504_ clknet_leaf_129_wb_clk_i team_02_WB.instance_to_wrap.top.DUT.read_data2\[7\]
+ _01378_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.dmmstore_co\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13716_ net1050 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
X_10928_ net383 _06356_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14696_ net1166 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16435_ clknet_leaf_90_wb_clk_i net1618 _01309_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.ru.imemaddr_co\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13647_ net1123 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16642__1213 vssd1 vssd1 vccd1 vccd1 _16642__1213/HI net1213 sky130_fd_sc_hd__conb_1
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10859_ net401 _06505_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16366_ clknet_leaf_102_wb_clk_i _02799_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.lcd.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_13578_ net1170 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15317_ clknet_leaf_115_wb_clk_i _01768_ _00275_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12772__A_N _05421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12529_ net1879 net351 net476 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16297_ clknet_leaf_97_wb_clk_i _02730_ _01240_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.a1.row2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16632__1380 vssd1 vssd1 vccd1 vccd1 net1380 _16632__1380/LO sky130_fd_sc_hd__conb_1
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15248_ clknet_leaf_34_wb_clk_i _01699_ _00206_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ clknet_leaf_22_wb_clk_i _01630_ _00137_ vssd1 vssd1 vccd1 vccd1 team_02_WB.instance_to_wrap.top.DUT.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10905__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout308 _06975_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_1
XANTENNA__09771__A2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout319 net322 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09740_ team_02_WB.instance_to_wrap.top.DUT.register\[6\]\[13\] net701 net632 team_02_WB.instance_to_wrap.top.DUT.register\[28\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10118__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

