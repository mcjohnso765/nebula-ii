* NGSPICE file created from team_02.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt team_02 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8]
+ gpio_in[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14]
+ gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20]
+ gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27]
+ gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XPHY_EDGE_ROW_176_Left_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ top.pad.keyCode\[5\] top.pad.keyCode\[4\] top.pad.keyCode\[6\] top.pad.keyCode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__or4b_1
X_06883_ top.DUT.register\[29\]\[25\] net787 net764 top.DUT.register\[19\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08622_ _03634_ _03724_ net291 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__mux2_1
XANTENNA__13840__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08553_ net320 _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nand2_1
XANTENNA__09287__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__B2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07298__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ top.DUT.register\[12\]\[14\] net647 net631 top.DUT.register\[27\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
X_08484_ net321 _02366_ _02449_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a21o_1
XANTENNA__07332__B _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07435_ _02551_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1071_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_185_Left_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout427_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07366_ top.DUT.register\[24\]\[5\] net586 net583 top.DUT.register\[4\]\[5\] _02482_
+ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06317_ top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] _01455_ top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__or4b_1
X_09105_ _04148_ _04149_ _04150_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07297_ top.DUT.register\[16\]\[1\] net724 net718 top.DUT.register\[9\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08163__B _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _04085_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06248_ net1357 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[6\] sky130_fd_sc_hd__and2_1
XFILLER_0_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 top.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net1 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XANTENNA__10913__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09546__Y _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 top.DUT.register\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 top.DUT.register\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07494__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold373 top.DUT.register\[11\]\[17\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 top.DUT.register\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 top.DUT.register\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 _04170_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_2
Xfanout831 net833 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12938__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _04622_ net360 net329 top.a1.dataIn\[28\] net364 vssd1 vssd1 vccd1 vccd1
+ _04924_ sky130_fd_sc_hd__a221o_1
Xfanout842 _01594_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout853 _04084_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_4
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_181_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout886 _01439_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_4
X_09869_ _04860_ _04861_ _04859_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout897 net899 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
Xhold1040 top.DUT.register\[9\]\[20\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1051 top.DUT.register\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ net125 net126 vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nand2_1
Xhold1062 top.DUT.register\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__C top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12880_ clknet_leaf_115_clk _00426_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1073 top.DUT.register\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 top.DUT.register\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 top.DUT.register\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07523__A _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ _05682_ _05686_ _05661_ _05666_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_197_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09278__A1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10220__Y _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ _05612_ _05614_ top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07828__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13501_ clknet_leaf_120_clk _01047_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ net1952 net154 net497 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ _05549_ _05551_ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ clknet_leaf_33_clk _00978_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ net167 net2146 net377 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ clknet_leaf_109_clk _00909_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10095__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ net181 net2186 net502 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12314_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] _01447_ top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a31o_1
XANTENNA__07461__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ clknet_leaf_95_clk _00840_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12245_ net1154 net612 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__nor2_1
XANTENNA__10823__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09202__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__Y _03473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07213__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _06007_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__xor2_2
XFILLER_0_208_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11127_ net924 net1295 net876 _05063_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a31o_1
X_11058_ net4 net862 net834 net1187 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__o22a_1
XFILLER_0_155_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08713__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net149 net1574 net450 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07433__A _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07819__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07220_ top.DUT.register\[13\]\[9\] net790 net802 top.DUT.register\[31\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08264__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07151_ top.DUT.register\[10\]\[12\] net726 net584 top.DUT.register\[24\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ _02112_ _02198_ net291 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07452__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10733__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07204__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout127 _05724_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_2
Xfanout138 _04208_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_2
Xfanout149 _04941_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
X_07984_ _03094_ _03096_ _03098_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09723_ net813 _04735_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__or2_2
X_06935_ top.DUT.register\[12\]\[22\] net735 net720 top.DUT.register\[26\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout377_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ net908 top.a1.state\[0\] top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04677_
+ sky130_fd_sc_hd__nor3b_1
X_06866_ net324 _01981_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__nand2_1
X_08605_ net477 _02662_ _02666_ net458 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__a22oi_1
X_06797_ top.DUT.register\[5\]\[30\] net603 net724 top.DUT.register\[16\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
X_09585_ net132 _04596_ _04612_ net917 vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout544_A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ net476 _02798_ _02799_ net458 _03632_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_193_Left_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10908__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _02833_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07418_ top.DUT.register\[3\]\[5\] net693 net662 top.DUT.register\[18\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
X_08398_ net273 _03508_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__or2_1
XANTENNA__07691__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ top.DUT.register\[16\]\[6\] net724 net762 top.DUT.register\[30\]\[6\] _02465_
+ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_150_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10360_ net1539 net249 net432 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06797__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ net330 net620 net1317 net887 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__a2bb2o_1
X_10291_ net1309 net265 net524 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__mux2_1
XANTENNA__10643__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ _05858_ _05864_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold170 top.DUT.register\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09735__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold192 top.ramaddr\[18\] vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 _01696_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_8
Xfanout672 net674 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_8
Xfanout683 _01670_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_4
XANTENNA__09499__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout694 _01664_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ clknet_leaf_29_clk _00478_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ clknet_leaf_32_clk _00409_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11058__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ _05631_ _05635_ _05637_ net129 vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__and4_1
XFILLER_0_201_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08636__X _03739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ clknet_leaf_20_clk _00340_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _05568_ _05598_ _05602_ _05603_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nor4_1
XFILLER_0_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10818__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _05520_ _05525_ _05519_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13415_ clknet_leaf_52_clk _00961_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10627_ net239 net2024 net376 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13346_ clknet_leaf_10_clk _00892_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09974__A2 _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10558_ net253 net1773 net503 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13277_ clknet_leaf_120_clk _00823_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ net264 net1917 net380 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__09187__B1 _04224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net1934 net867 net831 net127 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ _06013_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire345_A _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ top.DUT.register\[22\]\[3\] net554 net661 top.DUT.register\[18\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
XANTENNA__08259__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06651_ top.DUT.register\[1\]\[2\] net704 net624 top.DUT.register\[16\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XANTENNA__11049__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06582_ net746 _01653_ _01658_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__and3_4
X_09370_ net856 _01805_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08321_ _03332_ _03336_ net318 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10728__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _01736_ _01744_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__or2_1
XANTENNA__07673__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ _02313_ _02315_ _02317_ _02319_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08183_ net299 _02264_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06228__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ top.DUT.register\[10\]\[13\] net726 net750 top.DUT.register\[19\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XANTENNA__07425__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06779__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ top.DUT.register\[21\]\[16\] net608 net752 top.DUT.register\[17\]\[16\] _02181_
+ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a221o_1
XANTENNA__10463__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1034_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout494_A _04999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ top.DUT.register\[31\]\[18\] net667 net647 top.DUT.register\[12\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net919 net133 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06918_ top.DUT.register\[5\]\[23\] net600 net726 top.DUT.register\[10\]\[23\] _02034_
+ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a221o_1
X_07898_ top.DUT.register\[10\]\[24\] net646 net642 top.DUT.register\[9\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ net919 top.pc\[30\] _04661_ net911 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__o211a_1
X_06849_ top.DUT.register\[14\]\[26\] net794 net590 top.DUT.register\[20\]\[26\] _01965_
+ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06703__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ top.pc\[27\] _04583_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08519_ _02799_ _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10638__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09499_ net823 _04528_ _04531_ net132 net917 vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ _05363_ _05364_ _05346_ _05349_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _05313_ _05316_ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire347 _02304_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09405__B2 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ clknet_leaf_117_clk _00746_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xwire358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
X_10412_ net2277 net167 net516 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__mux2_1
XANTENNA__07416__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11392_ top.a1.dataIn\[27\] _05251_ top.a1.dataIn\[28\] vssd1 vssd1 vccd1 vccd1 _05253_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13131_ clknet_leaf_6_clk _00677_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10373__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ net1454 net181 net518 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10274_ net188 net2129 net434 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
X_13062_ clknet_leaf_21_clk _00608_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08916__A0 _03924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _05815_ _05842_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__or2_1
XANTENNA__12506__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 _05013_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06942__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_6
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input10_X net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ clknet_leaf_111_clk _00461_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08695__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12228__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ clknet_leaf_94_clk _00392_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09910__B _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10548__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ clknet_leaf_27_clk _00323_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09644__A1 _01920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08085__Y _03202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ top.a1.dataIn\[10\] _05579_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _05510_ _05512_ _05516_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_211_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold906 top.DUT.register\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 top.DUT.register\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold928 top.DUT.register\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ clknet_leaf_9_clk _00875_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10283__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 top.DUT.register\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09925__X _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08870_ _03030_ _03055_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nor2_1
XANTENNA__07186__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ top.DUT.register\[31\]\[28\] net669 _02937_ vssd1 vssd1 vccd1 vccd1 _02938_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06933__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07752_ top.DUT.register\[21\]\[31\] net571 net562 top.DUT.register\[20\]\[31\] _02868_
+ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a221o_1
XANTENNA__09006__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08135__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06703_ top.DUT.register\[6\]\[4\] net578 net693 top.DUT.register\[3\]\[4\] _01819_
+ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a221o_1
X_07683_ _02799_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__inv_2
X_09422_ _01595_ _02525_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nor2_1
XANTENNA__07894__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ _01630_ _01748_ _01750_ net400 net856 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09353_ _04392_ _04393_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nand2_1
XANTENNA__10458__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ _01661_ _01668_ _01674_ _01681_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__or4_1
XANTENNA__09635__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13565__RESET_B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08304_ _02845_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07646__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09284_ _02325_ _02775_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__xnor2_1
X_06496_ _01512_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__and2_2
XFILLER_0_28_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07110__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08235_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout507_A _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ _01740_ _03281_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07117_ top.DUT.register\[15\]\[14\] net805 net801 top.DUT.register\[31\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ top.DUT.register\[1\]\[22\] net704 net672 top.DUT.register\[19\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a22o_1
XANTENNA__08071__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ top.DUT.register\[14\]\[17\] net793 net585 top.DUT.register\[24\]\[17\] _02156_
+ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload90 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_12
XFILLER_0_140_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10921__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _01709_ net620 net1157 net888 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ net1510 net219 net481 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_206_Right_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__A1 _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ clknet_leaf_18_clk _00246_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06688__A1 top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ clknet_leaf_88_clk _01221_ net1015 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09776__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ net2241 net234 net408 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
X_12631_ clknet_leaf_112_clk _00177_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10368__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12562_ clknet_leaf_89_clk _00108_ net1016 vssd1 vssd1 vccd1 vccd1 top.pc\[27\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07101__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11513_ _05369_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ clknet_leaf_89_clk _00040_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11444_ _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07249__Y _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11375_ _05221_ _05228_ _05235_ top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1 _05236_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_189_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ clknet_leaf_14_clk _00660_ net987 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ net1531 net253 net519 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13045_ clknet_leaf_83_clk _00591_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_2__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10831__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ net258 net1981 net435 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07168__A2 _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ net263 net2063 net440 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06915__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07876__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ net1138 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07441__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10278__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ clknet_leaf_118_clk _00375_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06350_ _01461_ _01478_ _01479_ _01334_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__o22a_1
XFILLER_0_173_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06281_ top.ramload\[7\] net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08840__A2 _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08020_ top.DUT.register\[3\]\[19\] net691 net560 top.DUT.register\[20\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold703 top.DUT.register\[10\]\[23\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 top.DUT.register\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold736 top.DUT.register\[19\]\[28\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 top.DUT.register\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__A1 _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold758 top.DUT.register\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold769 top.DUT.register\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _04951_ _04952_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ _02979_ _03006_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__and2_1
XANTENNA__10741__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net269 _03791_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout192_A _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07804_ top.DUT.register\[21\]\[29\] net568 net671 top.DUT.register\[19\]\[29\] _02920_
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a221o_1
X_08784_ net903 top.pc\[21\] net538 _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07735_ _02366_ _02769_ _02692_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09856__A1 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07622__Y _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07666_ top.DUT.register\[4\]\[10\] net548 net659 top.DUT.register\[18\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08447__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ _04412_ _04426_ _04427_ _04425_ _02195_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a32o_1
X_06617_ _01388_ _01489_ _01722_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__o21a_1
XANTENNA__10188__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout624_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ _02704_ _02713_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07619__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ net854 _01748_ net619 _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_173_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06548_ top.DUT.register\[30\]\[0\] net696 net692 top.DUT.register\[3\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06479_ top.a1.instruction\[2\] _01514_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08218_ net298 _02132_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _04232_ _04235_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _01874_ _01877_ _02952_ _02929_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11160_ net55 net880 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ net156 net1874 net386 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
X_11091_ net1200 net879 net847 top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__a22o_1
XANTENNA__10651__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ net151 net1708 net530 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
Xhold30 top.a1.data\[0\] vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold52 top.a1.data\[9\] vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 net112 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold74 net124 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 _01192_ vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_69_clk _01326_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold96 _01166_ vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _05810_ _05820_ _05833_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or3b_1
XANTENNA__11103__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13732_ clknet_leaf_64_clk _01262_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_10__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09460__B net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ net1564 net156 net485 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XANTENNA__07858__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06429__X _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07322__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13663_ clknet_leaf_90_clk _01204_ net1003 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
X_10875_ net1449 net169 net492 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09887__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ clknet_leaf_21_clk _00160_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ clknet_leaf_55_clk _01135_ net1095 vssd1 vssd1 vccd1 vccd1 top.ramload\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12545_ clknet_leaf_98_clk _00091_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[10\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__09459__Y _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10826__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09023__A1_N _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ clknet_leaf_76_clk _00023_ net1082 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08035__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _05259_ net478 vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07389__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09783__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ top.a1.dataIn\[21\] top.a1.dataIn\[20\] top.a1.dataIn\[22\] vssd1 vssd1 vccd1
+ vccd1 _05219_ sky130_fd_sc_hd__o21a_1
XANTENNA__10561__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net1967 net182 net523 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__mux2_1
X_11289_ top.lcd.nextState\[1\] _01382_ _05141_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_169_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ clknet_leaf_31_clk _00574_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1050 net1073 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1073 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_177_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_206_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07561__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09838__A1 _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ _02627_ _02636_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__or2_2
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07313__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__A1 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07451_ top.DUT.register\[6\]\[6\] net578 net693 top.DUT.register\[3\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06402_ top.a1.instruction\[17\] net830 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__nand2_1
X_07382_ top.DUT.register\[28\]\[4\] net741 _01546_ top.DUT.register\[16\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a22o_1
X_09121_ _01600_ _04173_ _04172_ _04171_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__a211o_1
X_06333_ _01464_ _01465_ _01461_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o21a_1
XANTENNA__10736__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _03622_ _04104_ _03547_ _03579_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__and4b_1
X_06264_ net1192 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_170_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06515__A top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ top.DUT.register\[30\]\[21\] net696 net553 top.DUT.register\[22\]\[21\] _03119_
+ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08026__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 top.DUT.register\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
X_06195_ top.pc\[23\] vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
Xhold511 top.DUT.register\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 top.DUT.register\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold533 top.DUT.register\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09774__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 top.DUT.register\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 top.DUT.register\[4\]\[1\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__A1 _04941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 top.DUT.register\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top.DUT.register\[22\]\[15\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 top.DUT.register\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10471__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09954_ net818 _04640_ _04937_ net816 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ net461 _03982_ _03994_ net466 _03992_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ net816 _04874_ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a211o_1
Xhold1200 top.DUT.register\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1211 top.ramload\[18\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ net279 _02028_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09561__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08767_ net1395 net859 net836 _03863_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout741_A _01526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _02469_ _02587_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__nand2_1
XANTENNA__09280__B _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__Y _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08698_ _03208_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07304__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08501__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07649_ _02759_ _02761_ _02763_ _02765_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__or4_2
XFILLER_0_193_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ net239 net1800 net420 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09319_ _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08265__B1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_114_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10591_ net254 net2220 net424 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
X_12330_ top.lcd.cnt_500hz\[11\] _06122_ _06124_ net743 vssd1 vssd1 vccd1 vccd1 _01347_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08017__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ _06072_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11212_ top.a1.data\[4\] net796 _05030_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o21a_1
XANTENNA__11167__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__B1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12192_ _06035_ _06051_ _06050_ _06049_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08640__A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_11143_ net922 net1326 net874 _05071_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a31o_1
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__10381__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__B _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XANTENNA__06431__Y _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__07791__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
X_11074_ net21 net863 net835 net1285 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ net221 net2185 net529 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XANTENNA__08740__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13642__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _05802_ _05834_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__xor2_1
XANTENNA__08087__A _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13715_ clknet_leaf_66_clk _01245_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ net1805 net223 net485 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13646_ clknet_leaf_88_clk net1189 net1017 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
X_10858_ net1607 net239 net491 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08256__B1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13577_ clknet_leaf_64_clk _01118_ net1107 vssd1 vssd1 vccd1 vccd1 top.a1.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_105_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10556__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10789_ net254 net2258 net413 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ clknet_leaf_93_clk _00074_ net996 vssd1 vssd1 vccd1 vccd1 top.ramstore\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12459_ clknet_leaf_79_clk top.ru.next_FetchedInstr\[22\] net1085 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[22\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08559__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09646__A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10291__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
XANTENNA__09933__X _04920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _02066_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__nor2_4
XANTENNA__06990__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _04190_ _04679_ _04686_ net908 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__a22o_1
X_06882_ top.DUT.register\[6\]\[25\] net598 net774 top.DUT.register\[2\]\[25\] _01998_
+ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07534__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08621_ _03679_ _03723_ net313 vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08552_ _03303_ _03307_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07503_ top.DUT.register\[2\]\[14\] net683 net560 top.DUT.register\[20\]\[14\] _02619_
+ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08483_ _03590_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nor2_1
XANTENNA__08495__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_A _04923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07434_ net302 net342 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07365_ top.DUT.register\[29\]\[5\] net787 net598 top.DUT.register\[6\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a22o_1
XANTENNA__10466__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1064_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09104_ _01741_ _02879_ _04151_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09995__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06316_ top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\] top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__or4bb_1
XANTENNA__12902__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07296_ top.DUT.register\[12\]\[1\] net737 net603 top.DUT.register\[5\]\[1\] _02412_
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _04086_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__nand2_1
X_06247_ net1848 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[5\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07470__A1 _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09747__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 top.DUT.register\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold341 top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XANTENNA__08460__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold352 top.DUT.register\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 top.DUT.register\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 top.DUT.register\[27\]\[15\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 top.DUT.register\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 _01517_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
Xfanout832 net833 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_2
X_09937_ net154 net2138 net390 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_2
XANTENNA_fanout956_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _01614_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
Xfanout865 _05004_ vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_2
Xfanout887 net888 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_2
X_09868_ top.pc\[21\] _04511_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_2
Xhold1030 top.DUT.register\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 top.DUT.register\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 top.DUT.register\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03232_ _03894_ _03229_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08722__B2 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1063 top.DUT.register\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06733__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1074 top.DUT.register\[28\]\[6\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ top.pc\[14\] _04391_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1085 top.DUT.register\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ _05682_ _05686_ _05661_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a21oi_1
Xhold1096 top.DUT.register\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _05587_ _05588_ _05615_ _05619_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ clknet_leaf_16_clk _01046_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ net1766 net159 net498 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
X_11692_ net178 _05528_ _05540_ _05550_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__o32a_2
XFILLER_0_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3__f_clk_X clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13431_ clknet_leaf_112_clk _00977_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ net170 top.DUT.register\[21\]\[23\] net374 vssd1 vssd1 vccd1 vccd1 _00785_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10376__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08789__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13362_ clknet_leaf_107_clk _00908_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10574_ net183 net1594 net502 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12313_ net742 _06113_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13293_ clknet_leaf_115_clk _00839_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12244_ net1153 _06021_ net612 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ top.a1.dataIn\[2\] _06025_ _06031_ _06024_ vssd1 vssd1 vccd1 vccd1 _06036_
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08410__B1 _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06602__B _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11126_ net68 net883 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11057_ net3 net851 net850 net2232 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07516__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__A1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__A _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ net151 net1974 net452 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06724__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07433__B _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11959_ _05783_ _05815_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__and3b_1
XFILLER_0_175_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13629_ clknet_leaf_93_clk net1201 net995 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10286__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ top.DUT.register\[21\]\[12\] net608 net760 top.DUT.register\[30\]\[12\] _02266_
+ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _02155_ _02197_ net315 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07167__Y _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07608__B net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07755__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout128 _05724_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_1
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_14__f_clk_X clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ top.DUT.register\[15\]\[18\] net688 net623 top.DUT.register\[16\]\[18\] _03099_
+ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a221o_1
Xfanout139 net142 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06963__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net813 _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__nor2_1
X_06934_ top.DUT.register\[15\]\[22\] net805 net801 top.DUT.register\[31\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a22o_1
XANTENNA__13172__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07507__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__A _02305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ top.a1.halfData\[3\] _01385_ _01422_ top.a1.halfData\[5\] vssd1 vssd1 vccd1
+ vccd1 _04676_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_207_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06865_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10321__Y _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ net306 _03707_ _03699_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__a21oi_1
X_09584_ _04604_ _04610_ _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o21ai_1
X_06796_ top.DUT.register\[22\]\[30\] net606 net732 top.DUT.register\[23\]\[30\] _01912_
+ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08535_ _03640_ _03641_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ _02837_ _03546_ _02835_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ top.DUT.register\[28\]\[5\] net658 net645 top.DUT.register\[10\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10196__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ net301 _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout704_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09838__X _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07348_ top.DUT.register\[14\]\[6\] net794 net783 top.DUT.register\[3\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10924__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07279_ top.DUT.register\[21\]\[2\] net609 net593 top.DUT.register\[8\]\[2\] _02395_
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ net1298 net887 _03151_ net622 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__a22o_1
XANTENNA__07994__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ net1428 net258 net522 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold160 top.ramstore\[4\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 top.DUT.register\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 top.DUT.register\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 top.pad.button_control.r_counter\[12\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06954__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _01699_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_4
Xfanout651 net654 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
Xfanout662 _01690_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_8
Xfanout684 _01670_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ clknet_leaf_34_clk _00477_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06706__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ clknet_leaf_37_clk _00408_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11813_ _05669_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12793_ clknet_leaf_56_clk _00339_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11744_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06437__X _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07131__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11675_ _05520_ _05525_ _05519_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ clknet_leaf_45_clk _00960_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net245 net1651 net376 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13345_ clknet_leaf_44_clk _00891_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ net266 net2170 net503 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10834__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13830__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ clknet_leaf_101_clk _00822_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ net240 net1685 net379 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XANTENNA__13683__RESET_B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ net1480 net867 net833 _05761_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07198__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13612__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _06002_ _06005_ _06012_ _06003_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a22oi_2
XANTENNA__06945__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ net92 net878 net846 net1229 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_16_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12089_ _05937_ _05946_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__xor2_2
XANTENNA__07444__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08259__B _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06650_ top.DUT.register\[14\]\[2\] net664 net660 top.DUT.register\[18\]\[2\] _01766_
+ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07370__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06581_ net746 _01647_ _01658_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__and3_4
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ _03329_ _03347_ net284 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XANTENNA__07122__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08251_ _01736_ _01744_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_25_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07202_ top.DUT.register\[16\]\[10\] net723 net584 top.DUT.register\[24\]\[10\] _02318_
+ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ _03296_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07133_ top.DUT.register\[8\]\[13\] net592 net770 top.DUT.register\[27\]\[13\] _02249_
+ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a221o_1
XANTENNA__10744__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07976__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ top.DUT.register\[14\]\[16\] net792 net748 top.DUT.register\[1\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1027_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06936__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__inv_2
X_09705_ top.a1.halfData\[5\] _01480_ _04710_ net1102 vssd1 vssd1 vccd1 vccd1 _00120_
+ sky130_fd_sc_hd__o211a_1
X_06917_ top.DUT.register\[27\]\[23\] net770 net756 top.DUT.register\[3\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ top.DUT.register\[11\]\[24\] net702 net685 top.DUT.register\[2\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__a22o_1
XANTENNA__08169__B _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09636_ net134 _04651_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__o21ai_1
X_06848_ top.DUT.register\[12\]\[26\] net736 net774 top.DUT.register\[2\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07361__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07900__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ net918 top.pc\[26\] _04595_ net911 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06779_ top.DUT.register\[21\]\[29\] net608 net750 top.DUT.register\[19\]\[29\] _01883_
+ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10919__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ _02693_ _02772_ _03584_ _02692_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07113__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09498_ _04529_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_176_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ net309 _03557_ _03558_ _03554_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11460_ _05286_ _05302_ _05299_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__or3b_1
XANTENNA__08472__X _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
Xwire348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire359 _01897_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
X_10411_ net1845 net172 net513 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10654__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ top.a1.dataIn\[27\] top.a1.dataIn\[28\] _05251_ vssd1 vssd1 vccd1 vccd1 _05252_
+ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13130_ clknet_leaf_118_clk _00676_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07967__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ net2331 net183 net517 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
X_13061_ clknet_leaf_47_clk _00607_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_52_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ net194 net2101 net434 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ _05830_ _05844_ _05864_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or3_2
XANTENNA__06927__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_8
Xfanout492 _05000_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09341__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__B2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12914_ clknet_leaf_115_clk _00460_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12845_ clknet_leaf_113_clk _00391_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_61_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10829__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07711__B _02611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12776_ clknet_leaf_26_clk _00322_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ top.a1.dataIn\[10\] _05546_ _05579_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11658_ _05497_ _05514_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08823__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ net174 net2333 net423 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10564__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ _05413_ _05444_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07958__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold907 top.DUT.register\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ clknet_leaf_117_clk _00874_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold918 top.DUT.register\[4\]\[17\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 top.DUT.register\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_70_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13259_ clknet_leaf_3_clk _00805_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06918__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ top.DUT.register\[14\]\[28\] net665 net645 top.DUT.register\[10\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a22o_1
XANTENNA__09373__B _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ top.DUT.register\[26\]\[31\] net682 net657 top.DUT.register\[28\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08135__A2 _03251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ top.DUT.register\[8\]\[4\] net559 net661 top.DUT.register\[18\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a22o_1
XANTENNA__12746__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ _02797_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _04454_ _04457_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__xnor2_1
X_06633_ top.a1.instruction\[23\] _01634_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06697__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _02244_ _04391_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or2_1
X_06564_ top.DUT.register\[13\]\[0\] net676 net553 top.DUT.register\[22\]\[0\] _01678_
+ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08303_ _03279_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09283_ _04323_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06495_ top.a1.instruction\[0\] top.a1.instruction\[1\] top.a1.instruction\[2\] top.a1.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout235_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _01919_ net358 net325 vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08165_ _01739_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10474__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__B _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07116_ _02226_ _02228_ _02230_ _02232_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__or4_1
XANTENNA__07949__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08096_ top.DUT.register\[26\]\[22\] net680 net557 top.DUT.register\[8\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_12
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ top.DUT.register\[12\]\[17\] net735 net758 top.DUT.register\[2\]\[17\] _02163_
+ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a221o_1
Xclkload91 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_101_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__B1 _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06540__X _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net890 _01494_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_4
XANTENNA__07582__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ top.DUT.register\[26\]\[20\] net680 net639 top.DUT.register\[9\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09323__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ net1338 net226 net481 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07334__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07371__X _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09874__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ net357 _04643_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10891_ net1608 net238 net409 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
XANTENNA__10649__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ clknet_leaf_16_clk _00176_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ clknet_leaf_87_clk _00107_ net1018 vssd1 vssd1 vccd1 vccd1 top.pc\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11512_ _05333_ _05368_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ clknet_leaf_89_clk _00039_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08643__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11443_ top.a1.dataIn\[18\] net327 _05295_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10384__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06434__Y _01551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11374_ _05228_ _05230_ _05219_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_189_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ clknet_leaf_57_clk _00659_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10325_ net1829 net265 net520 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__mux2_1
X_13044_ clknet_leaf_98_clk _00590_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ net261 net2115 net436 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10187_ net243 net1863 net439 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08117__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11121__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07325__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07722__A _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ net1137 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_159_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07441__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ clknet_leaf_18_clk _00374_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08825__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12759_ clknet_leaf_112_clk _00305_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06280_ net1357 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[6\] sky130_fd_sc_hd__and2_1
XANTENNA__08553__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06625__X _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06851__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09936__X _04923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold704 top.DUT.register\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 top.DUT.register\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 top.DUT.register\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 top.DUT.register\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06603__A2 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _04951_ _04952_ _04192_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a21oi_1
Xhold748 top.DUT.register\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 top.DUT.register\[5\]\[26\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ net307 _03686_ _03571_ net395 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08852_ net274 _03943_ _03613_ net307 vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07564__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ top.DUT.register\[30\]\[29\] net695 net627 top.DUT.register\[29\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_108_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08783_ _03876_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__or3b_2
XFILLER_0_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08108__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07734_ _02612_ _02829_ _02850_ _02827_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a31o_1
XANTENNA__12109__A1_N top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07316__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09856__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07665_ top.DUT.register\[3\]\[10\] net691 net540 top.DUT.register\[5\]\[10\] _02781_
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a221o_1
XANTENNA__10469__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06616_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07596_ _02706_ _02708_ _02710_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__or4_2
XANTENNA__09608__A2 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _01595_ _01637_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06547_ net746 _01652_ _01656_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _02346_ _02668_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__nand2_1
XANTENNA__06682__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__A _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ top.a1.instruction\[6\] _01482_ top.a1.instruction\[2\] net914 vssd1 vssd1
+ vccd1 vccd1 _01595_ sky130_fd_sc_hd__nand4b_4
X_08217_ _03329_ _03332_ net317 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06842__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ _01808_ net337 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12203__A_N top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09993__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08148_ _03007_ _03263_ _03264_ _02958_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout986_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ top.DUT.register\[1\]\[17\] net704 net561 top.DUT.register\[20\]\[17\] _03195_
+ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a221o_1
XANTENNA__10932__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ net160 net1898 net388 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__mux2_1
X_11090_ net1214 net878 net846 top.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net156 net1643 net529 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
XANTENNA__07555__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 top.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top.a1.data\[3\] vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 top.a1.data\[8\] vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 net114 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net103 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_69_clk _01325_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold86 net94 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 top.DUT.register\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11992_ _05851_ _05852_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__or2_2
XANTENNA__07307__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__A2 _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13731_ clknet_leaf_66_clk _01261_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10943_ net1723 net159 net486 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XANTENNA__10379__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ net1926 net170 net489 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_13662_ clknet_leaf_90_clk _01203_ net1011 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ clknet_leaf_40_clk _00159_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13593_ clknet_leaf_54_clk _01134_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramload\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12544_ clknet_leaf_98_clk _00090_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[9\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06833__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ clknet_leaf_75_clk _00022_ net1082 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08035__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11426_ _05265_ _05278_ _05283_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__or4_1
XFILLER_0_151_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_6 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09783__A1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11357_ top.a1.dataIn\[0\] _04676_ net870 _05218_ vssd1 vssd1 vccd1 vccd1 _01274_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10842__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07717__A _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ net1628 net185 net522 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__mux2_1
X_11288_ top.a1.row2\[40\] _05157_ _05158_ top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1
+ _05159_ sky130_fd_sc_hd__a22o_1
XANTENNA__06621__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_33_clk _00573_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07436__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ net193 net2198 net382 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_206_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1058 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 net1064 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07010__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1073 net1121 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_2
XFILLER_0_174_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1084 net1091 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
Xfanout1095 net1111 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08548__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10289__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07450_ _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06401_ top.a1.instruction\[16\] net830 top.a1.instruction\[15\] vssd1 vssd1 vccd1
+ vccd1 _01518_ sky130_fd_sc_hd__and3b_2
XFILLER_0_201_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07381_ top.DUT.register\[21\]\[4\] net610 net749 top.DUT.register\[1\]\[4\] _02497_
+ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ top.a1.instruction\[13\] _01489_ _01610_ vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__a21oi_1
X_06332_ _01464_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09051_ _03456_ _03491_ _03519_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__and4_1
XFILLER_0_142_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06263_ top.ramload\[21\] net895 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ top.DUT.register\[1\]\[21\] net704 net680 top.DUT.register\[26\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold501 top.DUT.register\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_06194_ top.pc\[16\] vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
Xhold512 top.DUT.register\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top.DUT.register\[21\]\[31\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A1 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold534 top.DUT.register\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10752__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 top.DUT.register\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06802__Y _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold556 top.DUT.register\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold567 top.DUT.register\[16\]\[31\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 top.DUT.register\[21\]\[29\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold589 top.DUT.register\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _04643_ net361 net328 top.a1.dataIn\[29\] net363 vssd1 vssd1 vccd1 vccd1
+ _04938_ sky130_fd_sc_hd__a221o_1
XANTENNA__06531__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ _03009_ _03993_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_5_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _04525_ net360 net328 top.a1.dataIn\[22\] net363 vssd1 vssd1 vccd1 vccd1
+ _04876_ sky130_fd_sc_hd__a221o_1
XANTENNA__06250__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1201 top.DUT.register\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08835_ _02519_ _03902_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__or2_1
X_08766_ net902 top.pc\[20\] net538 _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07717_ _02469_ _02587_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nor2_1
XANTENNA__11097__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _03253_ _03777_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout734_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09988__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ top.DUT.register\[23\]\[8\] net566 net554 top.DUT.register\[22\]\[8\] _02764_
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10927__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ top.DUT.register\[15\]\[15\] net690 net649 top.DUT.register\[12\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09318_ _02284_ _04359_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or2_1
XANTENNA__07068__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ net268 net2016 net424 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _04293_ _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13600__Q top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06815__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12260_ top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] top.lcd.cnt_20ms\[2\] vssd1 vssd1
+ vccd1 vccd1 _06082_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09214__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11211_ _05026_ _05038_ net369 net404 net1244 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a32o_1
XANTENNA__09765__A1 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _06035_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07808__Y _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07776__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
X_11142_ net45 net881 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__and2_1
XANTENNA__07240__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
X_11073_ net20 net852 _05054_ net1456 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__a22o_1
XANTENNA__08999__A1_N _01709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__07528__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net226 net2151 net529 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07543__Y _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__B _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11088__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _05802_ _05834_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ clknet_leaf_63_clk _01244_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ net1520 net228 net487 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13645_ clknet_leaf_42_clk net1631 net1071 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
X_10857_ net2213 net246 net491 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__mux2_1
XANTENNA__10837__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13290__RESET_B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13576_ clknet_leaf_61_clk _01117_ net1107 vssd1 vssd1 vccd1 vccd1 top.a1.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10788_ net266 net2103 net412 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ clknet_leaf_84_clk _00073_ net1020 vssd1 vssd1 vccd1 vccd1 top.ramstore\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06806__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ clknet_leaf_79_clk top.ru.next_FetchedInstr\[21\] net1077 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__A2 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10572__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _01391_ net479 _05243_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a21bo_1
X_12389_ net1762 net920 net35 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_93_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07767__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06950_ _02051_ _02054_ _02057_ _02058_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06881_ top.DUT.register\[5\]\[25\] net603 net586 top.DUT.register\[24\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ net297 _02244_ _02265_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_124_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09381__B _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ net396 _02741_ _02742_ net476 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_178_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07502_ top.DUT.register\[29\]\[14\] net627 net623 top.DUT.register\[16\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07298__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ _02773_ net460 _03589_ net469 vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08495__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08495__B2 _03603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12491__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ _02479_ _02488_ _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__or3_4
XFILLER_0_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10747__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ top.DUT.register\[27\]\[5\] net772 _02480_ vssd1 vssd1 vccd1 vccd1 _02481_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ _04152_ _04153_ _04154_ _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__and4_1
X_06315_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[8\] _01449_ vssd1 vssd1 vccd1 vccd1
+ _01454_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07295_ top.DUT.register\[22\]\[1\] net606 net721 top.DUT.register\[26\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _01410_ _01778_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nand2_1
X_06246_ net1221 net895 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[4\] sky130_fd_sc_hd__and2_1
XFILLER_0_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09747__A1 _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10482__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 top.DUT.register\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
Xhold331 top.DUT.register\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07758__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08460__B net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 top.DUT.register\[28\]\[26\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 top.DUT.register\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top.DUT.register\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold375 top.DUT.register\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold386 top.DUT.register\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 _01554_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_4
XANTENNA_fanout684_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold397 top.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06430__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ _03995_ net454 net533 _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__o211a_4
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
Xfanout833 _05093_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_2
Xfanout855 _01614_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_2
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 _01440_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ top.pc\[21\] _04511_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__and2_1
Xhold1020 top.DUT.register\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_1
Xhold1031 top.DUT.register\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout899 _01435_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_2
Xhold1042 top.DUT.register\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11607__A top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1053 top.DUT.register\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net470 _03901_ _03905_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__a211o_1
XFILLER_0_169_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1064 top.DUT.register\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ top.pc\[13\] _04378_ _04790_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a21o_1
XANTENNA__07930__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 top.DUT.register\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 top.DUT.register\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 top.DUT.register\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ net398 _03844_ _03845_ _01730_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__o22ai_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _05589_ top.a1.dataIn\[9\] _05546_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__or3b_1
XANTENNA__07289__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ net2314 net163 net500 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11691_ _05501_ _05504_ _05528_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13430_ clknet_leaf_104_clk _00976_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10642_ net177 net2042 net375 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07446__C1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__A2 _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_8_clk _00907_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10573_ net189 net2295 net501 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07997__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ top.lcd.cnt_500hz\[5\] _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__xnor2_1
X_13292_ clknet_leaf_3_clk _00838_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07461__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08651__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__A1 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ net1164 _06032_ net612 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XANTENNA__10392__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12173__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06442__Y _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _06033_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08410__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07213__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08410__B2 _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06171__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__C_N _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net924 net1333 net877 _05062_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_166_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input33_X net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ net33 net862 net834 net1653 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__o22a_1
X_10007_ net154 net2020 net450 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07714__B _02611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07921__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07433__C _02549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _05740_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07730__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06488__B1 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ net2283 net164 net409 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10567__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11889_ _05748_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13628_ clknet_leaf_93_clk net1215 net995 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13559_ clknet_leaf_109_clk _01105_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07080_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07452__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07204__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout129 _05649_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
X_07982_ top.DUT.register\[30\]\[18\] net695 net639 top.DUT.register\[9\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a22o_1
X_06933_ top.DUT.register\[3\]\[22\] net782 net707 top.DUT.register\[7\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a22o_1
X_09721_ _01619_ _01627_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__nor2_1
XANTENNA__13559__RESET_B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ top.a1.halfData\[3\] net907 _01422_ top.a1.halfData\[5\] vssd1 vssd1 vccd1
+ vccd1 _04675_ sky130_fd_sc_hd__and4b_1
X_06864_ _01971_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__nor2_4
X_08603_ net283 _03513_ _03685_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _04604_ _04610_ net823 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a21oi_1
X_06795_ top.DUT.register\[3\]\[30\] net782 net765 top.DUT.register\[19\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout265_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08534_ _02800_ _03639_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XANTENNA__07911__Y _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ net469 _03559_ _03574_ net394 _03568_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a221o_1
XANTENNA__10477__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ top.DUT.register\[7\]\[5\] net575 net681 top.DUT.register\[26\]\[5\] _02532_
+ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ _03359_ _03507_ net290 vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06256__A top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07691__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10049__Y _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ top.DUT.register\[23\]\[6\] net732 net764 top.DUT.register\[19\]\[6\] _02463_
+ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07979__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ top.DUT.register\[2\]\[2\] net759 net757 top.DUT.register\[3\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
XANTENNA__06543__X _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09017_ net1256 net889 _03102_ net622 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__a22o_1
XANTENNA__06651__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06229_ top.ru.state\[4\] top.busy_o top.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 _01437_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__B _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09854__X _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 _01162_ vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _01165_ vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top.DUT.register\[15\]\[14\] vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 top.ramaddr\[19\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold194 top.ramaddr\[5\] vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10940__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _01703_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
Xfanout641 _01699_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_8
Xfanout652 net654 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
X_09919_ _04897_ _04899_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_148_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 net666 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_8
Xfanout674 _01683_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
Xfanout685 _01670_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout696 _01663_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_4
X_12930_ clknet_leaf_25_clk _00476_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07903__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_119_clk _00407_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _05653_ _05671_ _05637_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and3b_1
X_12792_ clknet_leaf_37_clk _00338_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _05598_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__or2_2
XFILLER_0_37_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ _05525_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13413_ clknet_leaf_45_clk _00959_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06890__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10625_ net249 net1754 net376 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13344_ clknet_leaf_12_clk _00890_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10556_ net258 net1568 net502 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06642__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13275_ clknet_leaf_0_clk _00821_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ net616 _04733_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nand2_1
XANTENNA__09187__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ net833 _05796_ _05797_ net868 net1193 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12157_ _05997_ _06007_ _06009_ _06014_ _06016_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__o32a_1
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11108_ net91 net882 net848 net1188 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XANTENNA__07725__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12088_ _05947_ _05948_ _05940_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08320__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ top.a1.data\[7\] net796 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__or2_1
XANTENNA__09895__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06580_ top.DUT.register\[17\]\[0\] net652 net648 top.DUT.register\[12\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a22o_1
XANTENNA__08556__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10297__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ _03279_ _03280_ _01739_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__or3b_1
XFILLER_0_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07673__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07201_ top.DUT.register\[23\]\[10\] net730 net707 top.DUT.register\[7\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06881__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08181_ net326 _02195_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13655__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ top.DUT.register\[23\]\[13\] net730 net756 top.DUT.register\[3\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09387__A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07425__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07063_ top.DUT.register\[24\]\[16\] net584 net758 top.DUT.register\[2\]\[16\] _02179_
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10760__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _03080_ _03081_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout382_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _04695_ _04702_ _04719_ _04720_ net1102 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__o311a_1
X_06916_ top.DUT.register\[14\]\[23\] net792 net748 top.DUT.register\[1\]\[23\] _02032_
+ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a221o_1
X_07896_ top.DUT.register\[6\]\[24\] net579 net689 top.DUT.register\[15\]\[24\] _03012_
+ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a221o_1
XANTENNA__09886__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net138 _04654_ _04658_ _04659_ net919 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__o221a_1
X_06847_ top.DUT.register\[8\]\[26\] net594 net582 top.DUT.register\[4\]\[26\] _01963_
+ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout647_A _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06778_ top.DUT.register\[7\]\[29\] net707 net756 top.DUT.register\[3\]\[29\] _01882_
+ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a221o_1
X_09566_ net137 _04588_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_195_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08517_ net1344 net858 net836 _03624_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ top.pc\[21\] _04484_ top.pc\[22\] vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10000__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net296 _01856_ _03460_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06872__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08379_ _03476_ _03482_ _03491_ net464 _03488_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__o221a_1
XANTENNA__10935__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire327 _05293_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire338 _02508_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10410_ net1389 net176 net514 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire349 _02283_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_116_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07416__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ top.a1.dataIn\[26\] _05231_ _05249_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__or3_1
XANTENNA__08613__B2 _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11609__A1_N top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10341_ net1718 net188 net517 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13060_ clknet_leaf_29_clk _00606_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ net195 net1905 net435 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12011_ _05856_ _05869_ _05871_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10670__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 _03370_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
XFILLER_0_205_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout471 _02516_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
Xfanout482 _05003_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_4
Xfanout493 _04999_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_6
X_12913_ clknet_leaf_9_clk _00459_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__Y _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12228__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ clknet_leaf_4_clk _00390_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12775_ clknet_leaf_49_clk _00321_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ top.a1.dataIn\[10\] _05579_ _05546_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__B2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11657_ net178 vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__inv_2
XANTENNA__10845__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_211_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ net181 net1938 net423 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__mux2_1
XANTENNA__06624__A _01733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _05443_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__nand2_1
Xhold908 top.DUT.register\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ clknet_leaf_23_clk _00873_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10539_ net193 net2162 net426 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__mux2_1
Xhold919 top.DUT.register\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ clknet_leaf_117_clk _00804_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06911__X _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09565__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _06059_ _06060_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10580__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ clknet_leaf_40_clk _00735_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07040__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ _02860_ _02862_ _02864_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__or4_1
X_06701_ _01811_ _01813_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__or3_1
X_07681_ _02325_ _02796_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_211_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08540__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ _04455_ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__and2b_1
X_06632_ top.a1.instruction\[10\] _01486_ net824 top.a1.instruction\[15\] vssd1 vssd1
+ vccd1 vccd1 _01749_ sky130_fd_sc_hd__a22o_1
XANTENNA__07894__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09351_ _02244_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nand2_1
X_06563_ net747 _01647_ _01649_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__and3_1
X_08302_ _01713_ _03280_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _04324_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nor2_1
XANTENNA__07646__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06494_ _01491_ _01610_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__nor2_1
XANTENNA__08843__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08233_ net293 _03348_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10755__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _03279_ _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__or2_2
XANTENNA__09548__C _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ top.DUT.register\[28\]\[14\] net738 net784 top.DUT.register\[29\]\[14\] _02231_
+ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a221o_1
X_08095_ top.DUT.register\[21\]\[22\] net569 net640 top.DUT.register\[9\]\[22\] _03211_
+ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08071__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload70 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_8
X_07046_ top.DUT.register\[13\]\[17\] net789 net767 top.DUT.register\[11\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
Xclkload81 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_8
Xclkload92 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout597_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ net891 _01494_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_145_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09308__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07948_ top.DUT.register\[13\]\[20\] net675 _03064_ vssd1 vssd1 vccd1 vccd1 _03065_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_199_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09580__A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ top.DUT.register\[8\]\[27\] net556 net667 top.DUT.register\[31\]\[27\] _02995_
+ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07812__B _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ _01898_ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__nand2_1
X_10890_ net1560 net244 net408 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _04577_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__and2_1
XANTENNA__13603__Q top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07098__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ clknet_leaf_87_clk _00106_ net1018 vssd1 vssd1 vccd1 vccd1 top.pc\[25\] sky130_fd_sc_hd__dfstp_1
XANTENNA__07637__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11511_ _05369_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__xor2_1
XANTENNA__10665__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_199_Left_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12491_ clknet_leaf_89_clk _00038_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ net327 _05295_ top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11373_ top.a1.dataIn\[24\] _05232_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_189_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13112_ clknet_leaf_33_clk _00658_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10324_ net2194 net258 net519 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_189_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13043_ clknet_leaf_96_clk _00589_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ net242 net2012 net435 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XANTENNA__06450__Y _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ net614 _04975_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_208_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07722__B _02549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ net1136 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__07876__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ clknet_leaf_0_clk _00373_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07089__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ clknet_leaf_105_clk _00304_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11709_ _05563_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__or2_1
XANTENNA__10575__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ clknet_leaf_10_clk _00235_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11260__A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 top.DUT.register\[26\]\[30\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_203_Left_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold716 top.DUT.register\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 top.DUT.register\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold738 top.DUT.register\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold749 top.DUT.register\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07800__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10148__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ net399 _02955_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__nor2_1
XANTENNA__09002__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ _03870_ _03942_ net294 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__mux2_1
X_07802_ top.DUT.register\[15\]\[29\] net687 net667 top.DUT.register\[31\]\[29\] _02918_
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a221o_1
X_08782_ net461 _03865_ _03867_ net465 vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_127_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07913__A _02023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _02563_ _02838_ _02588_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__or3b_1
XANTENNA__12967__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07664_ top.DUT.register\[31\]\[10\] net667 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06529__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ _04419_ _04420_ _04421_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06615_ _01721_ _01727_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nor2_2
X_07595_ top.DUT.register\[20\]\[15\] net562 net558 top.DUT.register\[8\]\[15\] _02711_
+ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ _04362_ _04364_ _04360_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__o21ai_1
X_06546_ net747 _01647_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__and3_4
XANTENNA__07619__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06827__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10485__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09265_ _02366_ _02748_ _04302_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o21ai_1
X_06477_ top.a1.instruction\[6\] _01482_ top.a1.instruction\[2\] net914 vssd1 vssd1
+ vccd1 vccd1 _01594_ sky130_fd_sc_hd__and4b_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08463__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _03330_ _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09196_ _04242_ _04245_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08147_ _01982_ _02978_ _03008_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__or3b_1
XANTENNA__08044__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08078_ top.DUT.register\[30\]\[17\] net696 net684 top.DUT.register\[2\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07029_ top.DUT.register\[21\]\[18\] net608 net584 top.DUT.register\[24\]\[18\] _02145_
+ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout979_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__B _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07004__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ net160 net2052 net530 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
Xhold10 top.a1.dataInTemp\[11\] vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 _01163_ vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 top.ramstore\[16\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 top.lcd.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold54 top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 net88 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _01169_ vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 _01190_ vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold98 top.a1.row1\[12\] vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _05783_ _05815_ _05819_ _05833_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__and4b_1
XFILLER_0_98_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13730_ clknet_leaf_66_clk _01260_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ net1562 net163 net488 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XANTENNA__07858__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ clknet_leaf_90_clk _01202_ net1011 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ net1832 net174 net490 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ clknet_leaf_28_clk _00158_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13592_ clknet_leaf_54_clk _01133_ net1096 vssd1 vssd1 vccd1 vccd1 top.ramload\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06818__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ clknet_leaf_81_clk _00089_ net1079 vssd1 vssd1 vccd1 vccd1 top.pc\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07491__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ clknet_leaf_76_clk _00021_ net1082 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06174__A top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _05256_ _05284_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__nand2_1
XANTENNA__08035__A2 _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07243__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ top.a1.row2\[0\] net868 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06461__X _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11079__X _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ net2300 net187 net521 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__mux2_1
XANTENNA__07717__B _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ top.lcd.nextState\[1\] top.lcd.nextState\[0\] _05152_ vssd1 vssd1 vccd1 vccd1
+ _05158_ sky130_fd_sc_hd__and3_1
XANTENNA__06621__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ clknet_leaf_12_clk _00572_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ net197 net1935 net383 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_206_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 net1050 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12412__Q top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1044 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_2
Xfanout1052 net1058 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_2
X_10169_ net1747 net191 net525 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1074 net1079 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08829__A _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1085 net1087 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1099 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ net72 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06400_ top.a1.instruction\[19\] net830 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ top.DUT.register\[12\]\[4\] net736 net762 top.DUT.register\[30\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06331_ _01333_ _01334_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__xor2_1
XANTENNA__06809__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ _01740_ _03364_ _03365_ _03419_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06262_ net1297 net895 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[20\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ top.DUT.register\[15\]\[21\] net688 net557 top.DUT.register\[8\]\[21\] _03117_
+ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a221o_1
XANTENNA__08026__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06193_ top.pc\[15\] vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
XANTENNA__09223__A1 _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 top.DUT.register\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold513 top.DUT.register\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 top.DUT.register\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07234__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09774__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 top.DUT.register\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 top.DUT.register\[17\]\[0\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 top.DUT.register\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 top.DUT.register\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 top.DUT.register\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _04933_ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ _02979_ _03963_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ net819 _04531_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1202 top.DUT.register\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net303 _03596_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout1002_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _03847_ _03855_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__or3b_2
XFILLER_0_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07716_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ net470 _03787_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06259__A top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ top.DUT.register\[19\]\[8\] net673 net653 top.DUT.register\[17\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07578_ _02690_ _02691_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06546__X _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ _02284_ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06529_ top.a1.instruction\[24\] net799 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09248_ top.pc\[8\] _02591_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_153_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08017__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ top.pc\[2\] top.pc\[3\] vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11210_ _05023_ _05036_ net369 net404 net1243 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a32o_1
X_12190_ _06044_ _06048_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09765__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_186_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net922 net1318 net874 _05070_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a31o_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
X_11072_ net19 net863 net835 net1324 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__o22a_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__clkbuf_4
X_10023_ net229 net2061 net530 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06751__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_201_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ clknet_leaf_62_clk _01243_ net1109 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[111\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_127_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10925_ net2312 net234 net487 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13644_ clknet_leaf_42_clk net1329 net1100 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
X_10856_ net2248 net251 net491 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13575_ clknet_leaf_61_clk _01116_ net1107 vssd1 vssd1 vccd1 vccd1 top.a1.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ net259 net2023 net412 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ clknet_leaf_89_clk _00072_ net1015 vssd1 vssd1 vccd1 vccd1 top.ramstore\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07464__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12407__Q top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10853__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ clknet_leaf_74_clk top.ru.next_FetchedInstr\[20\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[20\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07216__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11408_ _01391_ net479 vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12388_ _01403_ _06160_ net815 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ _05139_ _05150_ _05182_ net906 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06990__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13009_ clknet_leaf_10_clk _00555_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10523__A0 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ top.DUT.register\[16\]\[25\] net724 net583 top.DUT.register\[4\]\[25\] _01996_
+ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_145_Left_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ net828 _02615_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__nand2_2
X_08481_ net396 _02771_ _02770_ net476 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07432_ _02529_ _02548_ net827 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_4
XFILLER_0_9_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ top.DUT.register\[15\]\[5\] net807 net802 top.DUT.register\[31\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09102_ _03128_ _03154_ _03179_ _03205_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__and4_1
X_06314_ _01448_ _01450_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__or4_4
XANTENNA__07455__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ top.DUT.register\[18\]\[1\] net779 net594 top.DUT.register\[8\]\[1\] _02410_
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_198_Right_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06245_ net1902 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[3\] sky130_fd_sc_hd__and2_1
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09033_ _01410_ _01778_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__or2_1
XANTENNA__10763__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout308_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold310 top.DUT.register\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XANTENNA__09747__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 top.DUT.register\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 top.DUT.register\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 top.DUT.register\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 top.DUT.register\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 top.DUT.register\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top.DUT.register\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06261__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold387 top.DUT.register\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _01554_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
Xhold398 top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ net816 _04918_ _04919_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a31o_1
Xfanout812 _01516_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_2
Xfanout823 _01633_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 _05055_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_2
XANTENNA_fanout677_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _01453_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_2
XANTENNA__06981__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
X_09866_ top.pc\[20\] _04494_ _04853_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_181_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_2
Xhold1010 top.DUT.register\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 top.DUT.register\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07373__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net891 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_4
Xhold1032 top.DUT.register\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ _01746_ _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_163_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1043 top.DUT.register\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 top.DUT.register\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _04391_ net362 _04796_ _04769_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a211o_1
XANTENNA__06733__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__B _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 top.DUT.register\[27\]\[22\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 top.DUT.register\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09999__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10003__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _02109_ _03079_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__or2_1
XANTENNA__09004__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1098 top.DUT.register\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08679_ net466 _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__nor2_1
XANTENNA__10938__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10710_ net1663 net167 net499 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XANTENNA__07694__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _05532_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ net181 net2120 net376 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13360_ clknet_leaf_115_clk _00906_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_172_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10572_ net191 net1666 net501 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12311_ net742 _06111_ _06112_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10673__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ clknet_leaf_6_clk _00837_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09199__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ net1148 _06042_ net612 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ top.a1.dataIn\[2\] _06031_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11124_ net67 net884 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ net32 net851 net850 net2239 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_181_Left_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10006_ net161 net2321 net452 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06724__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ net125 net126 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10848__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net2189 net167 net408 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XANTENNA__07730__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07685__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ _05717_ net128 _05721_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13627_ clknet_leaf_75_clk net1228 net1084 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10839_ net1411 net181 net495 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_13558_ clknet_leaf_102_clk _01104_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ clknet_leaf_44_clk _00055_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10583__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13489_ clknet_leaf_9_clk _01035_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__A1 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06660__B2 top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08988__S _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ top.DUT.register\[21\]\[18\] net568 net683 top.DUT.register\[2\]\[18\] _03097_
+ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_130_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06963__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ net614 _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand2_4
X_06932_ net325 _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__or2_1
XANTENNA__08289__A _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__inv_2
X_06863_ _01975_ _01977_ _01979_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__or3_1
XANTENNA__07912__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ net306 _03705_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or2_1
X_09582_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06794_ top.DUT.register\[1\]\[30\] net780 _01910_ vssd1 vssd1 vccd1 vccd1 _01911_
+ sky130_fd_sc_hd__a21o_1
X_08533_ _02800_ _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__or2_1
XANTENNA__10758__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout160_A _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout258_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07676__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ net309 _03557_ _03573_ _03554_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07415_ top.DUT.register\[8\]\[5\] net558 net653 top.DUT.register\[17\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11162__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _03448_ _03506_ net315 vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XANTENNA__13431__Q top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_A _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07428__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ top.DUT.register\[29\]\[6\] net786 net774 top.DUT.register\[2\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10493__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ top.DUT.register\[13\]\[2\] net789 net727 top.DUT.register\[10\]\[2\] _02390_
+ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09016_ _03202_ net620 net1178 net887 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__a2bb2o_1
X_06228_ net905 _01436_ net34 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A _01529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 top.ramaddr\[2\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 top.DUT.register\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 top.ramaddr\[29\] vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 top.a1.row1\[9\] vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 top.a1.row1\[3\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 top.a1.row1\[109\] vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout961_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_2
Xfanout631 net634 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_4
XANTENNA__08936__A1_N _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06954__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout642 _01699_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_2
X_09918_ top.pc\[26\] _04590_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__xor2_1
Xfanout653 net654 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08199__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 net666 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
Xfanout686 _01670_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09849_ top.pc\[19\] _04477_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__or2_1
Xfanout697 _01663_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_198_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06706__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_leaf_17_clk _00406_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _05653_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nand2b_1
X_12791_ clknet_leaf_107_clk _00337_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10668__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11742_ _05555_ _05580_ _05567_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07667__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07131__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11673_ _05530_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ clknet_leaf_28_clk _00958_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07419__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net256 net1956 net376 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08662__A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__X _04163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ clknet_leaf_47_clk _00889_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10555_ net262 net2287 net504 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__mux2_1
XANTENNA__08092__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13274_ clknet_leaf_20_clk _00820_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10486_ net139 net1706 net507 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12225_ net1272 net867 net833 _05833_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07198__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _06014_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__or2_1
XFILLER_0_209_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08601__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06945__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ net90 net886 net849 net1630 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12087_ _05916_ _05921_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__nand2_1
X_11038_ net1218 _05048_ net480 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
XANTENNA__12420__Q top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09940__B _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07370__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07741__A _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_201_Right_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10578__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ clknet_leaf_119_clk _00535_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07122__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07200_ top.DUT.register\[5\]\[10\] net600 net580 top.DUT.register\[4\]\[10\] _02316_
+ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ net299 _02223_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07131_ top.DUT.register\[12\]\[13\] net734 net766 top.DUT.register\[11\]\[13\] _02247_
+ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06804__B _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07188__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ top.DUT.register\[22\]\[16\] net604 net766 top.DUT.register\[11\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
XANTENNA__09021__A1_N _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07830__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09583__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06936__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _02109_ _03079_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ top.a1.halfData\[3\] _01480_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__or2_1
X_06915_ top.DUT.register\[26\]\[23\] net719 net584 top.DUT.register\[24\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
X_07895_ top.DUT.register\[23\]\[24\] net566 net554 top.DUT.register\[22\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13709__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _04644_ _04646_ _04657_ net823 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a31o_1
XANTENNA__07897__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ top.DUT.register\[21\]\[26\] net609 net717 top.DUT.register\[9\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XANTENNA__08747__A _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net133 _04585_ _04592_ _04593_ net919 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o221a_1
XFILLER_0_179_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06777_ top.DUT.register\[29\]\[29\] net784 _01880_ _01893_ vssd1 vssd1 vccd1 vccd1
+ _01894_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout542_A _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ net902 top.pc\[9\] net537 _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09496_ top.pc\[21\] top.pc\[22\] _04484_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__and3_1
XANTENNA__08310__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07113__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08447_ net301 _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nor2_1
XANTENNA__06321__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09578__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08378_ _03489_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07329_ top.DUT.register\[21\]\[7\] net610 net772 top.DUT.register\[27\]\[7\] _02445_
+ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08074__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ net1555 net193 net518 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10951__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ net202 net1877 net434 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__mux2_1
X_12010_ _05853_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06927__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 _04961_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_6
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout472 _01746_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
XFILLER_0_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_8
Xfanout494 _04999_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
X_12912_ clknet_leaf_117_clk _00458_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_6_clk _00389_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10398__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_15__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ clknet_leaf_47_clk _00320_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06177__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06608__C _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ _05548_ _05579_ _05581_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11656_ _05511_ _05516_ _05512_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_37_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06464__X _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ net186 net1836 net422 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ _05444_ _05445_ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06624__B _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ clknet_leaf_110_clk _00872_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold909 top.DUT.register\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ net195 net2183 net427 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12415__Q top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10861__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ clknet_leaf_8_clk _00803_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10469_ net211 net1580 net506 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12208_ _06059_ _06062_ _06060_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a21oi_1
X_13188_ clknet_leaf_29_clk _00734_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06918__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _05975_ _05991_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__and2_1
XANTENNA_wire343_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06700_ top.DUT.register\[29\]\[4\] net629 _01814_ _01816_ vssd1 vssd1 vccd1 vccd1
+ _01817_ sky130_fd_sc_hd__a211o_1
X_07680_ _02325_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__and2_1
XANTENNA__07879__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07343__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__B2 _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ top.a1.instruction\[22\] _01634_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06551__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09350_ net854 _01750_ net619 _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__o22a_2
XANTENNA__13622__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10101__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ net746 _01653_ _01662_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__and3_1
X_08301_ _02845_ net460 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _02668_ top.pc\[10\] vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06493_ net912 top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__nor2_1
X_08232_ _03345_ _03347_ net317 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08056__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ net314 _02428_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07114_ top.DUT.register\[1\]\[14\] net781 net766 top.DUT.register\[11\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a22o_1
XANTENNA__07803__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08094_ top.DUT.register\[31\]\[22\] net668 net644 top.DUT.register\[10\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload60 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__10771__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ top.DUT.register\[22\]\[17\] net605 net731 top.DUT.register\[23\]\[17\] _02159_
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a221o_1
Xclkload71 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__clkinv_8
Xclkload82 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_fanout1032_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ net1364 net861 net839 _04081_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__a22o_1
XANTENNA__07582__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ top.DUT.register\[1\]\[20\] net703 net667 top.DUT.register\[31\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06790__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ top.DUT.register\[23\]\[27\] net564 net675 top.DUT.register\[13\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a22o_1
XANTENNA__06549__X _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07334__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09617_ _02613_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__nor2_4
X_06829_ top.DUT.register\[9\]\[27\] net715 net580 top.DUT.register\[4\]\[27\] _01945_
+ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a221o_1
XANTENNA__08196__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout924_A _01400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10011__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _01993_ _02002_ _04576_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or3_1
XFILLER_0_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10946__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09479_ _02090_ _04511_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11510_ _05285_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12490_ clknet_leaf_89_clk _00037_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08047__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ _05277_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_156_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ _05228_ _05230_ _01394_ _05220_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a211o_1
X_13111_ clknet_leaf_107_clk _00657_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10323_ net2193 net262 net520 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10681__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__B1 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ clknet_leaf_105_clk _00588_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ net614 _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__nand2_4
X_10185_ _04738_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_208_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11106__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _01857_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13284__RESET_B net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13645__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07325__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11121__A3 _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13875_ net1135 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06619__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12826_ clknet_leaf_15_clk _00372_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10856__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12757_ clknet_leaf_100_clk _00303_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08825__A2 top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06906__Y _02023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _05564_ _05565_ _05568_ _05524_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a211o_1
XFILLER_0_182_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ clknet_leaf_113_clk _00234_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _05497_ _05498_ top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_181_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08589__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold706 top.DUT.register\[14\]\[23\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 top.a1.row1\[15\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_120_clk _00855_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_96_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold728 top.DUT.register\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10591__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold739 top.DUT.register\[21\]\[3\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09002__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06370__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _03906_ _03941_ net317 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__mux2_1
X_07801_ top.DUT.register\[11\]\[29\] net699 net655 top.DUT.register\[28\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a22o_1
XANTENNA__07564__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ net311 net395 _03515_ _03873_ _01745_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a32o_1
XANTENNA__06772__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07732_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__inv_2
XANTENNA__07316__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07663_ top.DUT.register\[13\]\[10\] net675 net663 top.DUT.register\[14\]\[10\] _02779_
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ _04438_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_140_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06614_ _01712_ net475 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__or2_1
X_07594_ top.DUT.register\[22\]\[15\] net554 net625 top.DUT.register\[16\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
X_09333_ _04373_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ top.a1.instruction\[22\] top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01662_ sky130_fd_sc_hd__and2_2
XANTENNA__10766__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ top.pc\[9\] _04297_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__xnor2_1
X_06476_ net914 net913 _01485_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06545__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ net298 _02068_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__and2_1
XANTENNA__08029__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ _04242_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout505_A _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09777__B1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _03056_ _03262_ _02982_ _03009_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08077_ top.DUT.register\[7\]\[17\] net573 net644 top.DUT.register\[10\]\[17\] _03193_
+ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07028_ top.DUT.register\[26\]\[18\] net719 net766 top.DUT.register\[11\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13724__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 top.a1.data\[7\] vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 _01177_ vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 top.ramstore\[14\] vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _02881_ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 top.ramstore\[11\] vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold66 _01184_ vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net77 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _05815_ _05819_ _05833_ _05847_ _05817_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__a41oi_1
Xhold88 top.ramstore\[7\] vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold99 top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10941_ net1727 net166 net487 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ clknet_leaf_89_clk _01201_ net1015 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ net1487 net179 net490 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12611_ clknet_leaf_35_clk _00157_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08268__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ clknet_leaf_55_clk _01132_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramload\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10676__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12542_ clknet_leaf_80_clk _00088_ net1079 vssd1 vssd1 vccd1 vccd1 top.pc\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_148_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12473_ clknet_leaf_75_clk _00020_ net1084 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_49_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09768__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _05255_ _05279_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__xor2_1
XANTENNA_8 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11355_ net1150 net1115 net845 _05217_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__a31o_1
XANTENNA__08440__B1 _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10306_ net1910 net191 net521 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__mux2_1
XANTENNA__08991__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ top.lcd.nextState\[1\] top.lcd.nextState\[0\] _05141_ vssd1 vssd1 vccd1 vccd1
+ _05157_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13025_ clknet_leaf_45_clk _00571_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ net201 net1776 net382 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_2
Xfanout1031 net1034 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1044 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
Xfanout1053 net1058 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_58_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10168_ net1270 net196 net526 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA__06754__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1072 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1075 net1079 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1086 net1087 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_10099_ net206 net2212 net388 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13858_ net72 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ clknet_leaf_27_clk _00355_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_108_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13789_ clknet_leaf_70_clk _01314_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06330_ _01331_ _01332_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06261_ net2349 net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[19\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08000_ top.DUT.register\[18\]\[21\] net660 net628 top.DUT.register\[29\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__a22o_1
X_06192_ top.pc\[8\] vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold503 top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 top.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold525 top.DUT.register\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 top.DUT.register\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold547 top.DUT.register\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 top.DUT.register\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04934_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold569 top.DUT.register\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ net473 _03987_ _03991_ net471 _03990_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _04870_ _04872_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07537__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ net277 _03922_ _03925_ net270 _03770_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a32o_1
XFILLER_0_148_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1203 top.DUT.register\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout190_A _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout288_A _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ net461 _03841_ _03860_ net465 vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__o22a_1
X_07715_ _02830_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__or2_1
XANTENNA__11097__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ _03208_ net459 _03793_ net473 _03794_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout455_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06259__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ top.DUT.register\[2\]\[8\] net685 net649 top.DUT.register\[12\]\[8\] _02762_
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07170__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ _02693_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__inv_2
XANTENNA__10496__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_A _04082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09316_ net856 _01637_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06528_ top.a1.instruction\[24\] net799 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ _01413_ _02591_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06459_ top.DUT.register\[7\]\[0\] net708 net754 top.DUT.register\[18\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07658__X _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09178_ _04209_ _04221_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ top.DUT.register\[10\]\[16\] net643 net623 top.DUT.register\[16\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06722__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07776__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ net44 net880 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_101_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_11071_ net18 net852 _05054_ top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__a22o_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07528__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net234 net1616 net531 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _05804_ _05810_ _05813_ _05820_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__o41a_2
XFILLER_0_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13712_ clknet_leaf_63_clk _01242_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_10924_ net1714 net236 net487 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07161__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07700__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10855_ net2072 net254 net492 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__mux2_1
X_13643_ clknet_leaf_93_clk net1205 net996 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13574_ clknet_leaf_61_clk _01115_ net1107 vssd1 vssd1 vccd1 vccd1 top.a1.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ net263 net1765 net413 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__mux2_1
X_12525_ clknet_leaf_93_clk _00071_ net996 vssd1 vssd1 vccd1 vccd1 top.ramstore\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__Y _03772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13833__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12456_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[19\] net1085 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _05241_ net478 _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__o21ba_1
X_12387_ net815 _06159_ _06160_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07767__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11338_ net1222 net843 _05204_ net1114 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__o211a_1
XANTENNA__06975__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11269_ _05128_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ clknet_leaf_116_clk _00554_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06727__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11266__A top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07500_ net826 _02616_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__nor2_4
X_08480_ net305 _03588_ _03587_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07152__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07431_ _02538_ _02547_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__nor2_2
XFILLER_0_159_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07362_ _02472_ _02474_ _02476_ _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__or4_4
XFILLER_0_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08862__X _03954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ _02839_ _03231_ _03254_ _03279_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__and4_1
X_06313_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\] top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__or4b_1
XFILLER_0_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07293_ top.DUT.register\[27\]\[1\] net772 net764 top.DUT.register\[19\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a22o_1
X_09032_ _01409_ _01643_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__or2_1
X_06244_ net1947 net895 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[2\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 top.DUT.register\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold311 top.DUT.register\[15\]\[0\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06175_ top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_A _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold322 top.DUT.register\[30\]\[4\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold333 top.DUT.register\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 top.DUT.register\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13316__RESET_B net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold355 top.DUT.register\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 top.DUT.register\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold377 top.DUT.register\[15\]\[23\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 top.DUT.register\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _01554_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
XFILLER_0_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06430__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ net819 _04596_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_110_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold399 top.DUT.register\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 _01499_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_2
Xfanout824 _01616_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_2
Xfanout835 _05055_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_2
XANTENNA__07654__A _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ net184 net1673 net390 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__mux2_1
Xfanout857 _01613_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06718__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 top.DUT.register\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 _04681_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_181_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout572_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 _01439_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_2
Xhold1011 top.DUT.register\[10\]\[4\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 top.DUT.register\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 top.DUT.register\[5\]\[6\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _03565_ _03569_ _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07373__B _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1044 top.DUT.register\[18\]\[17\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net818 _04400_ _04766_ top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 _04796_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1055 top.DUT.register\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 top.DUT.register\[12\]\[5\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ _02109_ _03079_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 top.DUT.register\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1088 top.DUT.register\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 top.DUT.register\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout837_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand2_1
XANTENNA__07143__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07629_ net400 _01642_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10640_ net183 net1892 net374 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10954__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ net197 net2137 net502 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12310_ top.lcd.cnt_500hz\[4\] _01447_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07997__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ clknet_leaf_2_clk _00836_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ _06048_ net612 _06070_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10202__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ top.a1.dataIn\[2\] _06031_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06957__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net925 net1275 net877 _05061_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__Y _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ net31 net862 net834 net2226 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__o22a_1
XANTENNA__06709__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ net164 net2029 net453 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07382__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07570__Y _02687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ _05783_ _05807_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__o21a_1
XANTENNA__07134__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ net1471 net173 net406 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
X_11887_ _05716_ _05721_ net128 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or3b_1
XFILLER_0_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06627__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09778__X _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ net1825 net185 net494 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
X_13626_ clknet_leaf_88_clk net1220 net1016 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12418__Q top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10864__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13557_ clknet_leaf_83_clk _01103_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10769_ net197 net2060 net372 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12508_ clknet_leaf_88_clk _00054_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramstore\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13488_ clknet_leaf_116_clk _01034_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ clknet_leaf_54_clk top.ru.next_FetchedInstr\[2\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06948__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ top.DUT.register\[11\]\[18\] net699 net627 top.DUT.register\[29\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06931_ _02047_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09362__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ top.edg2.flip1 _01390_ _04190_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a21o_1
XANTENNA__10104__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ top.DUT.register\[26\]\[26\] net720 net776 top.DUT.register\[17\]\[26\] _01978_
+ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a221o_1
X_08601_ _03508_ _03704_ net283 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__mux2_1
XANTENNA__07912__A2 _03028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ net353 _04607_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nand2_1
X_06793_ top.DUT.register\[15\]\[30\] net806 net802 top.DUT.register\[31\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XANTENNA__09114__A1 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08532_ _03600_ _03638_ _02691_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08965__A2_N _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _01855_ net356 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout153_A _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ top.DUT.register\[23\]\[5\] net567 net546 top.DUT.register\[24\]\[5\] _02530_
+ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ _03312_ _03321_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07345_ top.DUT.register\[10\]\[6\] net729 net586 top.DUT.register\[24\]\[6\] _02461_
+ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout320_A _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09848__B _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06824__Y _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ top.DUT.register\[6\]\[2\] net597 net708 top.DUT.register\[7\]\[2\] _02392_
+ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a221o_1
X_09015_ _03251_ net621 net1171 net888 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06227_ top.ru.state\[2\] top.busy_o vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__and2_1
XANTENNA__06651__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold130 top.a1.row1\[120\] vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold141 top.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 top.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 top.a1.row1\[0\] vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A _01534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 net93 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold185 top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 top.DUT.register\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_6
Xfanout621 _04083_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_6
X_09917_ net163 top.DUT.register\[1\]\[25\] net393 vssd1 vssd1 vccd1 vccd1 _00147_
+ sky130_fd_sc_hd__mux2_1
Xfanout632 net634 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_4
Xfanout643 _01698_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_4
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 _01695_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
Xfanout676 net678 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10014__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout687 _01667_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_4
X_09848_ top.pc\[19\] _04477_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__nand2_1
Xfanout698 _01663_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07903__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ net220 net1647 net391 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _05635_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__xnor2_2
X_12790_ clknet_leaf_104_clk _00336_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11741_ _05554_ _05566_ _05568_ _05579_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_194_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11672_ _05532_ _05531_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and2b_1
XFILLER_0_165_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10623_ net268 net1878 net377 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
X_13411_ clknet_leaf_34_clk _00957_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10684__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06890__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08178__B1_N _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ clknet_leaf_37_clk _00888_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10554_ net242 net2339 net502 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ clknet_leaf_55_clk _00819_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06642__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ net143 net1671 net507 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ _05864_ _05094_ net867 net1239 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _05997_ _05999_ _06006_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__o31a_1
XANTENNA__09493__B _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11106_ net89 net886 net849 net1328 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a22o_1
X_12086_ _05909_ _05937_ _05945_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_88_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11037_ net864 _05046_ _05047_ net869 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1
+ _05048_ sky130_fd_sc_hd__a32o_1
XFILLER_0_204_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07355__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ clknet_leaf_16_clk _00534_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11939_ _05773_ _05785_ _05796_ _05797_ _05767_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a41o_1
XANTENNA__08855__B1 _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10594__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ clknet_leaf_79_clk _01150_ net1085 vssd1 vssd1 vccd1 vccd1 top.ramload\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06881__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07130_ top.DUT.register\[14\]\[13\] net792 net711 top.DUT.register\[25\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06373__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ top.DUT.register\[26\]\[16\] net719 net760 top.DUT.register\[30\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _02099_ _02108_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_79_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09702_ _04709_ _04714_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__or3b_1
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06914_ top.DUT.register\[22\]\[23\] net604 net596 top.DUT.register\[6\]\[23\] _02030_
+ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07894_ top.DUT.register\[24\]\[24\] net547 net543 top.DUT.register\[5\]\[24\] _03010_
+ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a221o_1
XANTENNA__12543__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07346__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06845_ net298 net354 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__nand2_1
X_09633_ _04644_ _04646_ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10769__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09564_ _04577_ _04580_ _04591_ net822 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a31o_1
X_06776_ top.DUT.register\[4\]\[29\] net580 net752 top.DUT.register\[17\]\[29\] _01892_
+ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08515_ net463 _03606_ _03622_ _03364_ _03620_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a221o_2
XFILLER_0_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _04526_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08846__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08446_ net287 _03434_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06321__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06872__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08377_ _02562_ _02846_ _03454_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__or3_1
XFILLER_0_190_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_A _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07328_ top.DUT.register\[17\]\[7\] net777 net762 top.DUT.register\[30\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07259_ top.DUT.register\[6\]\[3\] net599 net765 top.DUT.register\[19\]\[3\] _02375_
+ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_59_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10009__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10270_ net205 net1972 net436 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07585__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _04976_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_6
XANTENNA__08129__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _04961_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_21_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout462 _03368_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_8
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout484 _05003_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_4
Xfanout495 _04999_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_6
X_12911_ clknet_leaf_25_clk _00457_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_118_clk _00388_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12773_ clknet_leaf_39_clk _00319_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11724_ _05503_ _05547_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11655_ _05492_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09488__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ net188 net1992 net422 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
X_11586_ _05407_ _05440_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ clknet_leaf_114_clk _00871_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10537_ net199 net2203 net426 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10468_ net214 net1753 net505 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__mux2_1
X_13256_ clknet_leaf_24_clk _00802_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09565__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ net1808 net866 net831 _06066_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__a22o_1
X_13187_ clknet_leaf_35_clk _00733_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap333_A _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ net2211 net219 net514 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__mux2_1
X_12138_ _05965_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__xor2_4
XANTENNA__07040__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ _05881_ _05896_ _05899_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_193_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07328__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ top.a1.instruction\[9\] _01486_ net824 top.a1.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07471__B _02549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06561_ top.DUT.register\[26\]\[0\] net680 net557 top.DUT.register\[8\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ net472 net272 _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__or3_1
XANTENNA__10635__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ top.pc\[10\] _02668_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__nand2b_1
X_06492_ _01607_ _01608_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08231_ net298 _01981_ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08162_ net314 _02428_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09966__X _04950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07113_ top.DUT.register\[8\]\[14\] net592 net712 top.DUT.register\[25\]\[14\] _02229_
+ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ top.DUT.register\[15\]\[22\] net688 net632 top.DUT.register\[27\]\[22\] _03209_
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_6
X_07044_ top.DUT.register\[5\]\[17\] net601 net804 top.DUT.register\[15\]\[17\] _02160_
+ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a221o_1
XANTENNA__09005__B1 _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload72 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload72/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload83 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_12
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload94 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload94/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07567__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net905 top.pc\[31\] _03293_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout485_A _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ top.DUT.register\[8\]\[20\] net557 net549 top.DUT.register\[4\]\[20\] _03062_
+ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07877_ top.DUT.register\[15\]\[27\] net687 net548 top.DUT.register\[4\]\[27\] _02993_
+ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__a221o_1
XANTENNA__10499__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09616_ top.a1.instruction\[29\] net841 net618 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_178_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06828_ top.DUT.register\[27\]\[27\] net770 net748 top.DUT.register\[1\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09547_ _01993_ _02002_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__o21ai_1
X_06759_ top.DUT.register\[26\]\[28\] net721 _01861_ _01875_ vssd1 vssd1 vccd1 vccd1
+ _01876_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout917_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10626__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07098__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ _02090_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08429_ net472 net273 _03538_ _03371_ _02837_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload0 clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
X_11440_ net327 _05295_ _05274_ _05275_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10962__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__Y _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _05228_ _05230_ _05220_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_150_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ net1551 net240 net518 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__mux2_1
X_13110_ clknet_leaf_102_clk _00656_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07837__A _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ clknet_leaf_7_clk _00587_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09547__A1 _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _04959_ _04974_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nor2_2
XANTENNA__12465__RESET_B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ top.a1.instruction\[9\] top.a1.instruction\[10\] net744 vssd1 vssd1 vccd1
+ vccd1 _04974_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_100_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_208_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout270 _02202_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout281 net283 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
Xfanout292 _01774_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09116__X _04169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10202__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874_ net1134 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
X_12825_ clknet_leaf_44_clk _00371_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07089__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ clknet_leaf_97_clk _00302_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ _05523_ _05559_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__xor2_4
XFILLER_0_72_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12687_ clknet_leaf_19_clk _00233_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09786__X _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11638_ _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__A1 _03695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ _05375_ _05415_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07797__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 top.DUT.register\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 top.DUT.register\[9\]\[28\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_18_clk _00854_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07261__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold729 top.DUT.register\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ clknet_leaf_111_clk _00785_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07800_ top.DUT.register\[6\]\[29\] net576 net635 top.DUT.register\[25\]\[29\] _02916_
+ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a221o_1
X_08780_ _03875_ _03764_ _03874_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07731_ _02551_ _02558_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07662_ top.DUT.register\[9\]\[10\] net639 net631 top.DUT.register\[27\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a22o_1
XANTENNA__10112__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12494__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06613_ _01719_ _01728_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or2_1
X_09401_ top.pc\[17\] _04425_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_140_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07593_ top.DUT.register\[23\]\[15\] net566 net637 top.DUT.register\[25\]\[15\] _02709_
+ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08277__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06544_ top.DUT.register\[7\]\[0\] net573 net700 top.DUT.register\[11\]\[0\] _01655_
+ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a221o_1
X_09332_ _04353_ _04354_ _04355_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10619__Y _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ _04305_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_173_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06827__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06475_ net914 net913 _01485_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ net298 _02090_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nor2_1
X_09194_ _04243_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08145_ _02024_ _03029_ _03057_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__or3b_1
XANTENNA__09777__A1 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08076_ top.DUT.register\[5\]\[17\] net541 net652 top.DUT.register\[17\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07027_ top.DUT.register\[23\]\[18\] net730 net588 top.DUT.register\[20\]\[18\] _02143_
+ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a221o_1
XANTENNA__06460__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07004__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 top.pad.button_control.r_counter\[16\] vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 top.ramstore\[30\] vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 top.a1.data\[2\] vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08488__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ _02905_ _04044_ _01920_ _02901_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a2bb2o_1
Xhold45 top.ramstore\[12\] vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _01172_ vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 top.lcd.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ top.DUT.register\[1\]\[25\] net705 net634 top.DUT.register\[27\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a22o_1
Xhold78 _01174_ vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 _01168_ vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10940_ net2227 net171 net485 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XANTENNA__10022__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_203_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ net1335 net183 net489 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08494__Y _03603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ clknet_leaf_12_clk _00156_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13590_ clknet_leaf_55_clk _01131_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramload\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ clknet_leaf_83_clk _00087_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06818__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6__f_clk_X clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07491__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ clknet_leaf_89_clk _00019_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11423_ _05255_ _05279_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10692__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07779__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11354_ net845 _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07243__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10305_ net1512 net197 net523 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__mux2_1
X_11285_ top.a1.row1\[0\] _05154_ _05155_ top.a1.row1\[16\] vssd1 vssd1 vccd1 vccd1
+ _05156_ sky130_fd_sc_hd__a22o_1
X_13024_ clknet_leaf_13_clk _00570_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09782__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ net204 net1867 net384 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
Xfanout1010 net1014 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net39 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_4
Xfanout1032 net1034 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
X_10167_ net1509 net201 net525 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_2
Xfanout1054 net1058 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_2
Xfanout1065 net1067 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_4
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
X_10098_ net209 net1599 net386 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
Xfanout1087 net1089 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_2
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07703__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13857_ net72 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10867__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ clknet_leaf_25_clk _00354_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ clknet_leaf_70_clk _01313_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11271__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06809__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12739_ clknet_leaf_35_clk _00285_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06260_ net2350 net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
XFILLER_0_199_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07482__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06191_ top.pc\[6\] vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold504 top.DUT.register\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 top.DUT.register\[23\]\[10\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07234__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 top.DUT.register\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold537 top.DUT.register\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09082__C_N _03888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold548 top.DUT.register\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09950_ top.pc\[29\] _04643_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_1
Xhold559 top.DUT.register\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10107__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ net307 _03654_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__nor2_1
X_09881_ _04870_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11727__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ net286 _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__or2_1
Xhold1204 top.DUT.register\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08763_ _03858_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout183_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ _02448_ _02611_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08694_ net398 _03205_ _03204_ net477 vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07940__A _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10777__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ top.DUT.register\[31\]\[8\] net669 net625 top.DUT.register\[16\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ _02346_ _02689_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ net841 _01635_ net619 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__a21oi_1
X_06527_ _01486_ _01600_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09246_ top.pc\[7\] _02567_ _04283_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a21o_1
X_06458_ net811 _01527_ net808 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__and3_2
XFILLER_0_133_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09177_ _04086_ _04089_ _04226_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__a21o_1
X_06389_ top.pad.button_control.r_counter\[16\] top.pad.button_control.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__nand2_1
XANTENNA__13635__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08128_ top.DUT.register\[4\]\[16\] net548 net544 top.DUT.register\[24\]\[16\] _03244_
+ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07225__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06291__A top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ _03169_ _03171_ _03173_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or4_1
XANTENNA__10017__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__09806__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
X_11070_ net17 net863 net835 net1241 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__o22a_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net236 top.DUT.register\[3\]\[7\] net531 vssd1 vssd1 vccd1 vccd1 _00193_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09922__A1 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09107__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__A _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11972_ _05823_ _05827_ _05828_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__a21o_2
X_13711_ clknet_leaf_63_clk _01241_ net1106 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ net2323 net246 net488 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__mux2_1
XANTENNA__10687__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_197_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13642_ clknet_leaf_89_clk net1823 net1013 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
X_10854_ net1737 net265 net492 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ clknet_leaf_61_clk top.a1.nextHex\[4\] net1110 vssd1 vssd1 vccd1 vccd1 _01381_
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ net243 net1973 net411 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12524_ clknet_leaf_93_clk _00070_ net995 vssd1 vssd1 vccd1 vccd1 top.ramstore\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07464__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06672__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12455_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[18\] net1074 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ top.a1.dataIn\[21\] _05244_ _05245_ net479 vssd1 vssd1 vccd1 vccd1 _05267_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07216__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ top.pad.button_control.r_counter\[15\] _06157_ vssd1 vssd1 vccd1 vccd1 _06160_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08719__A1_N net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11337_ top.a1.row1\[108\] _05183_ _05192_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13686__RESET_B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ net900 net906 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09913__A1 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ clknet_leaf_21_clk _00553_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10219_ _04732_ _04974_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nor2_2
X_11199_ net870 net865 _05095_ _05102_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__or4_1
XFILLER_0_206_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10597__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07430_ _02540_ _02542_ _02544_ _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ top.DUT.register\[21\]\[5\] net611 net764 top.DUT.register\[19\]\[5\] _02477_
+ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08101__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06312_ top.lcd.cnt_500hz\[8\] top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] top.lcd.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__or4b_1
X_09100_ _02741_ _02771_ _02822_ _03054_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07292_ net297 net342 _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07455__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ net918 _01386_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__or2_1
XANTENNA__06663__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06243_ net1759 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[1\] sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09974__X _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06174_ top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09601__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold312 top.DUT.register\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold323 top.ramaddr\[3\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 top.DUT.register\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold345 top.a1.row1\[1\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 top.DUT.register\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top.DUT.register\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold378 top.DUT.register\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07494__X _02611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 top.DUT.register\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _04606_ net360 net328 top.a1.dataIn\[27\] net363 vssd1 vssd1 vccd1 vccd1
+ _04920_ sky130_fd_sc_hd__a221o_1
Xfanout803 _01554_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_4
Xfanout814 _06133_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_209_Left_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout825 net827 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout398_A _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09904__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07654__B _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout847 net848 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_2
X_09864_ _03862_ net454 net533 _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__o211a_2
Xfanout858 net860 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_2
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 top.DUT.register\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 top.DUT.register\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08815_ net269 _03751_ _03908_ net278 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__a22o_1
XANTENNA__11176__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 top.DUT.register\[18\]\[18\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ net214 net1606 net390 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
Xhold1034 top.DUT.register\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 top.DUT.register\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 top.DUT.register\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 top.DUT.register\[29\]\[5\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net310 _03473_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__and2_1
Xhold1078 top.DUT.register\[26\]\[10\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 top.DUT.register\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
X_08677_ _03257_ _03776_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _02743_ _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__nand2_2
XANTENNA__10300__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07694__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12920__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ top.DUT.register\[23\]\[9\] net566 net629 top.DUT.register\[29\]\[9\] _02675_
+ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10570_ net201 net2077 net501 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06573__X _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06654__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ top.pc\[6\] top.pc\[7\] _04254_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ net1147 net612 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12171_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11122_ net66 net884 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and2_1
Xhold890 top.DUT.register\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_166_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11053_ net30 net862 net834 net1357 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__o22a_1
XANTENNA__07906__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ net167 net1918 net453 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_199_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _05781_ _05807_ _05782_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12198__A top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06908__B _02023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10210__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10906_ net1363 net176 net407 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07685__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11886_ _05745_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nand2_1
X_13625_ clknet_leaf_59_clk net1235 net1071 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06893__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ top.DUT.register\[27\]\[19\] net187 net493 vssd1 vssd1 vccd1 vccd1 _00973_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06483__X _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13556_ clknet_leaf_97_clk _01102_ net1003 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10768_ net201 net1903 net370 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09831__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06645__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ clknet_leaf_76_clk _00053_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramstore\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07739__B _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ clknet_leaf_20_clk _01033_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ net1922 net215 net497 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09794__X _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12438_ clknet_leaf_54_clk top.ru.next_FetchedInstr\[1\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10880__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12369_ net1748 _06146_ _06148_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06930__Y _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire366_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06930_ _02042_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__nor2_4
X_06861_ top.DUT.register\[23\]\[26\] net731 net712 top.DUT.register\[25\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
X_08600_ _03611_ _03703_ net295 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__mux2_1
X_06792_ _01902_ _01904_ _01906_ _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__or4_4
X_09580_ net353 _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__or2_1
XANTENNA__09114__A2 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08531_ _02690_ _02770_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10120__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ _03570_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__nand2_1
XANTENNA__07676__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07413_ top.DUT.register\[6\]\[5\] net578 net641 top.DUT.register\[9\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06884__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ net309 _03504_ _03500_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_34_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout146_A _04950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ top.DUT.register\[1\]\[6\] net780 net714 top.DUT.register\[25\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07428__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07275_ top.DUT.register\[12\]\[2\] net735 net767 top.DUT.register\[11\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ _02714_ net621 net1155 net890 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__a2bb2o_1
X_06226_ net895 top.ru.next_dready net34 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__or3b_1
XFILLER_0_14_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09586__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 top.DUT.register\[7\]\[17\] vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 top.ramaddr\[22\] vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 top.DUT.register\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 top.ramaddr\[25\] vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08260__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 _01189_ vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 top.ramstore\[13\] vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
Xhold197 top.ramaddr\[16\] vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 _01522_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_4
XFILLER_0_186_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09916_ net535 _04896_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__and3_2
Xfanout622 _04082_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_6
Xfanout644 _01698_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout666 _01686_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_8
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_8
X_09847_ top.pc\[18\] _04460_ _04839_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 _01667_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
Xfanout699 _01660_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09778_ _03669_ net454 net533 _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_161_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08729_ _03361_ _03449_ net304 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11740_ _05524_ _05560_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10030__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07667__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__X _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06875__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _05472_ _05526_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10965__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13410_ clknet_leaf_10_clk _00956_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ net257 net2017 net375 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__07419__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ clknet_leaf_118_clk _00887_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10553_ net616 _04962_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__nand2_1
XANTENNA__08092__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13272_ clknet_leaf_38_clk _00818_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10484_ net149 net1769 net505 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ net1519 net868 net832 _05895_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__a22o_1
XANTENNA__07575__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ _05988_ _05995_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__xnor2_1
X_11105_ net1204 net879 net847 top.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 _01184_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10205__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ _05909_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nor2_1
XANTENNA_input31_X net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ top.a1.dataInTemp\[10\] net798 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ clknet_leaf_0_clk _00533_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ _05772_ _05785_ _05796_ _05797_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__nand4_4
XFILLER_0_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10875__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ _05703_ net127 _05705_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a21o_1
XANTENNA__09949__B _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09301__Y _04345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ clknet_leaf_79_clk _01149_ net1085 vssd1 vssd1 vccd1 vccd1 top.ramload\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08607__A1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__B2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ clknet_leaf_33_clk _01085_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08083__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07060_ top.DUT.register\[15\]\[16\] net804 net800 top.DUT.register\[31\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07830__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12720__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ net828 _03078_ net468 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__o21a_1
XANTENNA__10115__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _04696_ _04698_ _04703_ _04692_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__o22a_1
X_06913_ top.DUT.register\[13\]\[23\] net788 net707 top.DUT.register\[7\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
X_07893_ top.DUT.register\[13\]\[24\] net677 net650 top.DUT.register\[12\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09632_ _01919_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__xor2_1
X_06844_ _01953_ _01956_ _01958_ _01960_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__nor4_1
XANTENNA__07897__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _04577_ _04580_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a21oi_1
X_06775_ top.DUT.register\[8\]\[29\] net592 net584 top.DUT.register\[24\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08514_ _02695_ _03621_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__xnor2_1
X_09494_ _04509_ _04513_ _04512_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06857__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net293 _03438_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout430_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _02846_ _03454_ _02562_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06609__B1 _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ top.DUT.register\[13\]\[7\] net790 net721 top.DUT.register\[26\]\[7\] _02443_
+ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09271__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08074__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__B2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07282__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ top.DUT.register\[13\]\[3\] net790 net778 top.DUT.register\[18\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07821__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06209_ _01423_ _01428_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07189_ net323 _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09023__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06570__Y _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_8
Xfanout441 _04976_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 _04961_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _03367_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
Xfanout474 _01745_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
Xfanout485 _05002_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_8
Xfanout496 _04999_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
X_12910_ clknet_leaf_93_clk _00456_ net998 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12841_ clknet_leaf_28_clk _00387_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_169_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08837__A1 _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12772_ clknet_leaf_28_clk _00318_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11723_ _05543_ _05581_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06848__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10695__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11654_ _05495_ _05513_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ net192 net1772 net422 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11585_ _05444_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ clknet_leaf_115_clk _00870_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07273__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ net204 net1943 net428 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13255_ clknet_leaf_53_clk _00801_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_178_Left_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net216 net1888 net505 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__mux2_1
XANTENNA__09014__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12206_ _06058_ _06064_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07025__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13186_ clknet_leaf_12_clk _00732_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ net1828 net223 net513 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__mux2_1
X_12137_ top.a1.dataIn\[3\] _05981_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12068_ _05901_ _05924_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_205_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11019_ net1167 _05034_ net480 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
XANTENNA__07879__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06551__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06560_ _01659_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__nor2_4
XANTENNA__08864__A _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06491_ net913 _01599_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08230_ net324 _02003_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ _03265_ _03267_ _03270_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__nand4_1
XFILLER_0_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ top.DUT.register\[6\]\[14\] net596 net580 top.DUT.register\[4\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a22o_1
XANTENNA__11060__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07264__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ top.DUT.register\[3\]\[22\] net692 net652 top.DUT.register\[17\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a22o_1
XANTENNA__07803__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload40 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_8
X_07043_ top.DUT.register\[6\]\[17\] net597 net581 top.DUT.register\[4\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload51 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_6
Xclkload62 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload62/X sky130_fd_sc_hd__clkbuf_8
Xclkload73 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09005__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_16
Xclkload95 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_12
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ _04061_ _04078_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ top.DUT.register\[7\]\[20\] net572 net687 top.DUT.register\[15\]\[20\] _03061_
+ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08516__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06790__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ top.DUT.register\[1\]\[27\] net703 net699 top.DUT.register\[11\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a22o_1
XANTENNA__08110__Y _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ net134 _04640_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__nor2_1
X_06827_ top.DUT.register\[15\]\[27\] net804 net800 top.DUT.register\[31\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout645_A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ net840 _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_4
X_06758_ top.DUT.register\[6\]\[28\] net598 net594 top.DUT.register\[8\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09477_ net618 _04510_ _02614_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_191_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08428_ net396 _02834_ _02835_ net475 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_6
XANTENNA__13552__RESET_B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ net293 _01943_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09244__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11051__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07255__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06581__X _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ net617 _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__nor2_4
XFILLER_0_143_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07837__B _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06741__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07007__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ clknet_leaf_116_clk _00586_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09547__A2 _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10252_ net140 net2282 net384 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__mux2_1
XANTENNA__08014__A _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13855__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ top.a1.instruction\[9\] top.a1.instruction\[10\] net744 vssd1 vssd1 vccd1
+ vccd1 _04973_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_208_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 _04747_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11106__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _02203_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_2
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13873_ net1133 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12824_ clknet_leaf_33_clk _00370_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12755_ clknet_leaf_110_clk _00301_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06475__Y _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11706_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12686_ clknet_leaf_93_clk _00232_ net998 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11637_ _05456_ _05463_ _05491_ _05459_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a22o_2
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07246__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09786__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13222__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06932__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11568_ _05372_ _05427_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13307_ clknet_leaf_0_clk _00853_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold708 top.DUT.register\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ net140 net1767 net380 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__mux2_1
Xhold719 top.DUT.register\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ _05320_ _05322_ _05328_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a21oi_1
X_13238_ clknet_leaf_102_clk _00784_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ clknet_leaf_8_clk _00715_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07763__A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06772__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ net281 net343 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07661_ top.DUT.register\[11\]\[10\] net699 net568 top.DUT.register\[21\]\[10\] _02777_
+ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ top.pc\[17\] _04425_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06612_ _01719_ _01728_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_140_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ top.DUT.register\[30\]\[15\] net697 net629 top.DUT.register\[29\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _04371_ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06543_ net746 _01656_ _01658_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__and3_4
XFILLER_0_192_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07485__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09262_ _04306_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06474_ _01584_ _01588_ _01589_ _01590_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__nor4_1
XANTENNA__09772__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ _03327_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08029__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ top.pc\[4\] _01833_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10916__X _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07938__A _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _02068_ _03228_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09777__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__B2 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08075_ _03185_ _03187_ _03189_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07026_ top.DUT.register\[17\]\[18\] net752 net750 top.DUT.register\[19\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout595_A _01551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 _01369_ vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net1996 net861 net839 _04063_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__a22o_1
Xhold24 _01191_ vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net122 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 _01173_ vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07928_ top.DUT.register\[20\]\[25\] net563 net551 top.DUT.register\[4\]\[25\] _03044_
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a221o_1
XANTENNA__10303__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 net123 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold79 top.a1.data\[10\] vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10847__A1 _04941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _02969_ _02971_ _02973_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ net2131 net189 net489 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09529_ _04558_ _04559_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_158_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08268__A2 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07476__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ clknet_leaf_80_clk _00086_ net1079 vssd1 vssd1 vccd1 vccd1 top.pc\[5\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_80_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12471_ clknet_leaf_59_clk _00018_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.debounce
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10973__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08976__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ _05165_ _05184_ _05210_ net1114 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__or4b_1
XFILLER_0_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10304_ net2156 net199 net521 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11284_ _05133_ _05153_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nor2_1
X_13023_ clknet_leaf_23_clk _00569_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ net211 net1634 net382 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
XANTENNA__09782__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08679__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 net1002 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
Xfanout1011 net1014 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_2
Xfanout1022 net1023 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
X_10166_ net1245 net205 net527 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XANTENNA__06754__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1050 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_2
Xfanout1055 net1057 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
Xfanout1077 net1078 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_2
XANTENNA__10213__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10097_ net214 net2109 net387 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
Xfanout1099 net1111 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07703__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13856_ net72 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ clknet_leaf_44_clk _00353_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09303__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ clknet_leaf_71_clk _01312_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ top.a1.halfData\[1\] _05005_ _05018_ net865 vssd1 vssd1 vccd1 vccd1 _05019_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12738_ clknet_leaf_15_clk _00284_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07467__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ clknet_leaf_120_clk _00215_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07219__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06190_ top.pc\[3\] vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold505 top.DUT.register\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 top.DUT.register\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__A2 _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 top.DUT.register\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 top.DUT.register\[4\]\[3\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold549 top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
X_08900_ net279 _02518_ _03439_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__a31o_1
X_09880_ _04860_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _03884_ _03923_ net318 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__mux2_1
Xhold1205 top.DUT.register\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06745__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ _03083_ _03857_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__nand2_1
XANTENNA__08876__X _03967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ _02448_ _02611_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nor2_1
X_08693_ net304 _03362_ _03792_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout176_A _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ top.DUT.register\[1\]\[8\] net705 net570 top.DUT.register\[21\]\[8\] _02760_
+ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07170__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07432__S net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07575_ _02346_ _02689_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__and2_1
XANTENNA__09447__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09314_ _04353_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06526_ _01613_ _01642_ _01639_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_75_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09245_ net918 top.pc\[7\] _04292_ top.testpc.en_latched vssd1 vssd1 vccd1 vccd1
+ _00088_ sky130_fd_sc_hd__o211a_1
X_06457_ top.DUT.register\[25\]\[0\] net712 net758 top.DUT.register\[2\]\[0\] _01573_
+ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a221o_1
XANTENNA__09867__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout510_A _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08263__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _04086_ _04089_ _04226_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__a21oi_1
X_06388_ _01502_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ top.DUT.register\[19\]\[16\] net671 net635 top.DUT.register\[25\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06291__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08058_ top.DUT.register\[7\]\[23\] net573 net691 top.DUT.register\[3\]\[23\] _03174_
+ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06984__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ top.DUT.register\[13\]\[19\] net788 net723 top.DUT.register\[16\]\[19\] _02125_
+ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a221o_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_101_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10020_ net244 net2345 net531 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ top.a1.dataIn\[2\] top.a1.dataIn\[0\] top.a1.dataIn\[1\] vssd1 vssd1 vccd1
+ vccd1 _05832_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ clknet_leaf_63_clk _01240_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net2001 net251 net488 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07697__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ clknet_leaf_89_clk net1233 net1015 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10853_ net1355 net259 net491 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13572_ clknet_leaf_61_clk top.a1.nextHex\[3\] net1110 vssd1 vssd1 vccd1 vccd1 _01380_
+ sky130_fd_sc_hd__dfrtp_1
X_10784_ net616 _04979_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nand2_4
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ clknet_leaf_90_clk _00069_ net1003 vssd1 vssd1 vccd1 vccd1 top.ramstore\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12454_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[17\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ _05245_ net479 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__nand2_2
X_12385_ top.pad.button_control.r_counter\[15\] _06157_ vssd1 vssd1 vccd1 vccd1 _06159_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10208__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11336_ top.a1.row1\[60\] _05140_ _05188_ top.a1.row2\[12\] _05202_ vssd1 vssd1 vccd1
+ vccd1 _05203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06975__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ _05131_ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08177__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ clknet_leaf_92_clk _00552_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08177__B2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ net140 net2270 net440 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_105_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11198_ net1614 _05102_ _05096_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
XANTENNA__06727__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10149_ net141 net2095 net444 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09732__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13655__RESET_B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10878__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13839_ clknet_leaf_42_clk _01362_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09429__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ top.DUT.register\[16\]\[5\] _01545_ net777 top.DUT.register\[17\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_114_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06311_ top.lcd.cnt_500hz\[11\] _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07291_ net321 net339 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ net1287 net887 _02877_ net622 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__a22o_1
X_06242_ net1210 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[0\] sky130_fd_sc_hd__and2_1
XFILLER_0_127_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10118__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06173_ top.a1.dataIn\[24\] vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XANTENNA__12537__RESET_B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold302 top.DUT.register\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 top.DUT.register\[28\]\[31\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 top.DUT.register\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold335 top.DUT.register\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 top.DUT.register\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 top.DUT.register\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _04914_ _04915_ _04917_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__or3_1
Xhold368 top.DUT.register\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 top.DUT.register\[8\]\[8\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout804 _01553_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
Xfanout815 _06133_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout826 net827 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_8
X_09863_ _04171_ _04486_ _04855_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a211o_1
Xfanout837 net839 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_2
XANTENNA__08112__A _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA__06718__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_181_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _03825_ _03907_ net293 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
Xhold1002 top.DUT.register\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 top.DUT.register\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 top.DUT.register\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _03715_ net454 net533 _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__o211a_2
Xhold1035 top.DUT.register\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 top.DUT.register\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 top.DUT.register\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net303 _03473_ _03475_ _03571_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o31a_1
XFILLER_0_197_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10788__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 top.DUT.register\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 top.DUT.register\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout558_A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _03257_ _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_200_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07627_ net346 _02740_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_132_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_A _01545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07558_ top.DUT.register\[3\]\[9\] net693 net681 top.DUT.register\[26\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06509_ _01598_ _01623_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__nand2_1
XANTENNA__09597__B _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ top.DUT.register\[24\]\[7\] net546 net637 top.DUT.register\[25\]\[7\] _02605_
+ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _01412_ net853 net873 _04276_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_106_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10028__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _01778_ _02428_ _04210_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06406__A1 top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _06023_ _06026_ _06028_ _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_141_Left_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06957__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ net925 net1462 _01440_ _05060_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a31o_1
Xhold880 top.DUT.register\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold891 top.DUT.register\[26\]\[8\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_166_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ net29 net851 net850 net1848 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__a22o_1
XANTENNA__06709__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ net170 net2332 net450 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10698__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06590__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11954_ _05806_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_150_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08331__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08331__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ net1370 net179 net407 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ _05735_ _05739_ _05737_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08882__A2 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13624_ clknet_leaf_42_clk net1300 net1071 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
X_10836_ net1286 net192 net494 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XANTENNA__09788__A top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13555_ clknet_leaf_110_clk _01101_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08095__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10767_ net204 net1811 net372 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12506_ clknet_leaf_75_clk _00052_ net1084 vssd1 vssd1 vccd1 vccd1 top.ramstore\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07842__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13486_ clknet_leaf_95_clk _01032_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ net1611 net218 net497 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
X_12437_ clknet_leaf_54_clk top.ru.next_FetchedInstr\[0\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ top.pad.button_control.r_counter\[9\] _06146_ net814 vssd1 vssd1 vccd1 vccd1
+ _06148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_196_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06948__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11319_ net906 _05150_ _05186_ _05185_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12299_ net1142 _06105_ net1118 vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_130_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06860_ top.DUT.register\[16\]\[26\] net725 net761 top.DUT.register\[30\]\[26\] _01976_
+ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06791_ top.DUT.register\[8\]\[30\] net594 net777 top.DUT.register\[17\]\[30\] _01907_
+ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a221o_1
XANTENNA__06658__Y _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ net304 _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10401__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08461_ net307 net356 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__nand2_2
XFILLER_0_159_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07412_ top.a1.instruction\[26\] net854 _02527_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_159_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08392_ net301 _03503_ _03502_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12789__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07343_ top.DUT.register\[17\]\[6\] net777 _02459_ vssd1 vssd1 vccd1 vccd1 _02460_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08086__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07274_ top.DUT.register\[15\]\[2\] net804 net800 top.DUT.register\[31\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
X_09013_ net1183 net889 _02637_ net622 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06225_ top.busy_o top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 top.ru.next_iready sky130_fd_sc_hd__and2b_1
XFILLER_0_170_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 top.a1.row1\[104\] vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 top.ru.state\[4\] vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold132 top.busy_o vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 top.DUT.register\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold154 top.ramaddr\[7\] vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 top.ramaddr\[21\] vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 top.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08113__Y _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 top.ramaddr\[14\] vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 net603 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_8
Xfanout612 net613 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_4
Xhold198 top.ramaddr\[0\] vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11187__B _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09915_ net817 _04900_ _04901_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a31o_1
Xfanout623 net626 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_8
Xfanout634 _01702_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09889__A1 _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _01698_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout656 net658 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_8
Xfanout667 net668 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
X_09846_ net193 net1923 net391 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__mux2_1
XANTENNA__08010__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 _01679_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_4
XANTENNA__07364__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07681__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ top.a1.dataIn\[11\] _04766_ _04769_ _04779_ vssd1 vssd1 vccd1 vccd1 _04780_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ top.DUT.register\[29\]\[20\] net785 net727 top.DUT.register\[10\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout842_A _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ _03750_ _03825_ net295 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
XANTENNA__10311__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08659_ _02718_ _03740_ _02719_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _05479_ _05521_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06584__X _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ net262 net2292 net376 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09895__X _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ clknet_leaf_16_clk _00886_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10552_ net140 net2069 net428 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__mux2_1
XANTENNA__13858__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ clknet_leaf_111_clk _00817_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ _04932_ top.DUT.register\[16\]\[28\] net508 vssd1 vssd1 vccd1 vccd1 _00630_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12222_ net2276 net868 net832 _05924_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__a22o_1
X_12153_ _06002_ _06006_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ net87 net882 net848 net1822 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a22o_1
X_12084_ _05940_ _05941_ _05934_ _05938_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a211o_1
X_11035_ top.a1.data\[6\] net797 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2_1
XANTENNA__08001__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_X net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10221__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12986_ clknet_leaf_14_clk _00532_ net987 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13869__1129 vssd1 vssd1 vccd1 vccd1 _13869__1129/HI net1129 sky130_fd_sc_hd__conb_1
X_11937_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11868_ _05703_ _05705_ net127 vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09311__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net1652 net263 net496 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13607_ clknet_leaf_54_clk _01148_ net1077 vssd1 vssd1 vccd1 vccd1 top.ramload\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08068__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ _05627_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09804__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13538_ clknet_leaf_11_clk _01084_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10891__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ clknet_leaf_120_clk _01015_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ top.DUT.register\[5\]\[20\] net540 _03063_ _03068_ _03077_ vssd1 vssd1 vccd1
+ vccd1 _03078_ sky130_fd_sc_hd__a2111oi_1
X_09700_ top.a1.halfData\[2\] _01480_ _04717_ net1102 vssd1 vssd1 vccd1 vccd1 _00118_
+ sky130_fd_sc_hd__o211a_1
X_06912_ top.DUT.register\[15\]\[23\] net804 net801 top.DUT.register\[31\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
X_07892_ _03007_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__nand2_4
XANTENNA__07346__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ _02613_ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nor2_2
XFILLER_0_207_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06843_ top.DUT.register\[26\]\[27\] net719 net584 top.DUT.register\[24\]\[27\] _01959_
+ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a221o_1
XANTENNA__10131__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _01981_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__xor2_1
X_06774_ _01885_ _01886_ _01888_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_143_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08513_ _02770_ _03600_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__and2b_1
XFILLER_0_188_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09493_ _02068_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__xor2_1
XFILLER_0_203_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout256_A _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08444_ _02203_ _03552_ _03553_ net274 vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08375_ net472 net273 _03485_ _03486_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout423_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07326_ top.DUT.register\[1\]\[7\] net781 net732 top.DUT.register\[23\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a22o_1
XANTENNA__07806__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ top.DUT.register\[5\]\[3\] net602 net722 top.DUT.register\[26\]\[3\] _02373_
+ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06208_ top.a1.halfData\[5\] net920 _01421_ _01426_ vssd1 vssd1 vccd1 vccd1 _01428_
+ sky130_fd_sc_hd__or4_2
XFILLER_0_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07188_ net346 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout792_A _01529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1120_X net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08782__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06793__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _04994_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_6
Xfanout431 net433 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_6
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_8
Xfanout453 _04961_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 net467 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_4
XANTENNA__06579__X _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 _01730_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 _05002_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09731__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_8
X_09829_ top.pc\[17\] _04445_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__nand2_1
XANTENNA__08300__A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10041__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_26_clk _00386_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12771_ clknet_leaf_30_clk _00317_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10976__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11722_ _05543_ _05581_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ _05495_ _05513_ _05492_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10604_ net195 net2143 net423 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ _05408_ _05434_ _05410_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_6_clk _00869_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10535_ net208 net1729 net426 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06761__Y _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ clknet_leaf_48_clk _00800_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08034__X _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10466_ net220 net2316 net505 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12205_ net1436 net866 net831 _06065_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ clknet_leaf_43_clk _00731_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10216__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10397_ net1385 net231 net515 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
X_12136_ _05995_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2_2
XANTENNA__09970__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06784__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _05876_ _05925_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07328__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net864 _05032_ _05033_ net869 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1
+ _05034_ sky130_fd_sc_hd__a32o_1
XFILLER_0_204_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07989__A_N _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09740__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10886__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ clknet_leaf_27_clk _00515_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08864__B _03954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06490_ top.a1.instruction\[12\] _01601_ _01488_ vssd1 vssd1 vccd1 vccd1 _01607_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ _03181_ _03274_ _03275_ _03276_ _03060_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a41o_1
XFILLER_0_83_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07111_ top.DUT.register\[12\]\[14\] net735 net725 top.DUT.register\[16\]\[14\] _02227_
+ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _03204_ _03205_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload30 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload41 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_2
X_07042_ top.DUT.register\[8\]\[17\] net593 net708 top.DUT.register\[7\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
Xclkload52 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__09005__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload63 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinv_4
Xclkload74 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload85 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_2_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload96 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_8
XANTENNA__10126__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__inv_2
XANTENNA__06775__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07944_ top.DUT.register\[30\]\[20\] net695 net655 top.DUT.register\[28\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08516__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08516__B2 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _02985_ _02987_ _02989_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__or4_1
XFILLER_0_207_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout373_A _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ net284 _01942_ _01900_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a21o_1
X_09614_ _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_178_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09545_ top.a1.instruction\[25\] net842 net618 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10796__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06757_ _01869_ _01871_ _01872_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout638_A _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _01595_ _01642_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ top.a1.instruction\[16\] net824 _01804_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_191_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ _03413_ _03537_ net289 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_2
XANTENNA__08144__A_N _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout805_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06294__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ net301 _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__nor2_1
Xclkload2 clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09101__D _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07309_ top.DUT.register\[11\]\[1\] net769 net586 top.DUT.register\[24\]\[1\] _02425_
+ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08289_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_210_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10320_ top.a1.instruction\[7\] top.a1.instruction\[8\] _04181_ net744 vssd1 vssd1
+ vccd1 vccd1 _04982_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_104_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13868__1128 vssd1 vssd1 vccd1 vccd1 _13868__1128/HI net1128 sky130_fd_sc_hd__conb_1
X_10251_ net144 net2107 net385 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10036__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07558__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net1951 net141 net527 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XANTENNA__06766__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout250 _04756_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_208_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net264 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
Xfanout283 _01855_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net296 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
X_13872_ net1132 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_159_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07191__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12823_ clknet_leaf_111_clk _00369_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ clknet_leaf_105_clk _00300_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ _05564_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__and2_1
XANTENNA__07494__A1 _02610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ clknet_leaf_113_clk _00231_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13836__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11636_ _05481_ _05489_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a21o_2
XFILLER_0_112_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11567_ _05427_ _05372_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07797__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ net143 net2199 net380 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__mux2_1
X_13306_ clknet_leaf_15_clk _00852_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 top.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ _05322_ _05328_ _05330_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__and3_2
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ clknet_leaf_81_clk _00783_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10449_ net1483 net154 net509 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ clknet_leaf_116_clk _00714_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _05962_ _05979_ _05950_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__mux2_1
X_13099_ clknet_leaf_6_clk _00645_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire341_A _02407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ top.DUT.register\[8\]\[10\] net556 net635 top.DUT.register\[25\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a22o_1
XANTENNA__07182__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06611_ _01720_ _01727_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07591_ top.DUT.register\[21\]\[15\] net570 net645 top.DUT.register\[10\]\[15\] _02707_
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10069__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ top.pc\[13\] _04359_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06542_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09261_ _02748_ top.pc\[9\] vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__and2b_1
X_06473_ top.DUT.register\[22\]\[0\] net605 net767 top.DUT.register\[11\]\[0\] _01572_
+ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_173_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ net298 _02048_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nor2_1
X_09192_ top.pc\[4\] _01833_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__nor2_1
XANTENNA__06682__X _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _03207_ _03255_ _03206_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout219_A _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08074_ top.DUT.register\[14\]\[17\] net664 net549 top.DUT.register\[4\]\[17\] _03190_
+ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a221o_1
XANTENNA__06996__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__A _03229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ top.DUT.register\[22\]\[18\] net604 net756 top.DUT.register\[3\]\[18\] _02139_
+ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06460__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1030_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06748__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 top.a1.dataInTemp\[9\] vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _04061_ _04062_ net905 top.pc\[30\] vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__a2bb2o_1
Xhold25 top.a1.dataInTemp\[8\] vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top.lcd.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ top.DUT.register\[15\]\[25\] net690 net658 top.DUT.register\[28\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__a22o_1
Xhold58 top.ramload\[12\] vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 top.a1.data\[11\] vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06289__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ top.DUT.register\[11\]\[26\] net701 net570 top.DUT.register\[21\]\[26\] _02974_
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a221o_1
XANTENNA__07173__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06809_ top.DUT.register\[1\]\[31\] net780 net777 top.DUT.register\[17\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _02905_ _02881_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout922_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06920__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _02024_ _04557_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_158_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ net840 _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__nor2_2
XFILLER_0_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12470_ clknet_leaf_74_clk top.ru.next_read_i net1088 vssd1 vssd1 vccd1 vccd1 top.Ren
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11421_ _05280_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07779__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11352_ net1255 net843 _05215_ net1114 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06987__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10303_ net1460 net203 net523 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13866__A top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283_ _05137_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_18_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13022_ clknet_leaf_32_clk _00568_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10234_ net212 net2145 net382 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XANTENNA__07864__A _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_2
Xfanout1012 net1014 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10165_ net1349 net209 net525 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
Xfanout1023 net1030 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_210_Right_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1034 net1050 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_2
Xfanout1045 net1047 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_2
XANTENNA__07951__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1067 net1072 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
X_10096_ net218 net1597 net386 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1089 net1090 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07164__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__A2 _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13855_ net72 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ clknet_leaf_19_clk _00352_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09303__B _04345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10998_ top.a1.dataInTemp\[1\] net798 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__or2_1
X_13786_ clknet_leaf_65_clk _01311_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12737_ clknet_leaf_44_clk _00283_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ clknet_leaf_16_clk _00214_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11619_ _05473_ _05477_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nor3_1
XFILLER_0_182_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ clknet_leaf_111_clk _00145_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08967__B2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 top.DUT.register\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06978__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold517 top.DUT.register\[6\]\[0\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12453__Q top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 top.DUT.register\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 top.DUT.register\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08719__B2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _02025_ _02049_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__nand2_1
XANTENNA__10404__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1206 top.DUT.register\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ _03083_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__or2_1
X_07712_ _02468_ _02587_ _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nand3_1
X_08692_ net269 _03612_ _03791_ net278 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a22o_1
XANTENNA__07155__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07643_ top.DUT.register\[30\]\[8\] net697 net677 top.DUT.register\[13\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a22o_1
XANTENNA__06902__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout169_A _04895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07574_ _02346_ _02688_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__and2_1
X_13867__1127 vssd1 vssd1 vccd1 vccd1 _13867__1127/HI net1127 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_24_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09313_ _04354_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__and2b_1
X_06525_ top.a1.instruction\[21\] net824 _01641_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_196_Left_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ net133 _04279_ _04291_ net918 vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_62_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06456_ top.DUT.register\[27\]\[0\] net771 net761 top.DUT.register\[30\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _04086_ _04089_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__and3_1
X_06387_ top.pad.button_control.r_counter\[8\] _01504_ top.pad.button_control.r_counter\[10\]
+ top.pad.button_control.r_counter\[9\] vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_153_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ top.DUT.register\[9\]\[16\] net639 net627 top.DUT.register\[29\]\[16\] _03242_
+ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06969__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ top.DUT.register\[5\]\[23\] net541 net627 top.DUT.register\[29\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_186_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09001__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ top.DUT.register\[18\]\[19\] net754 net748 top.DUT.register\[1\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_168_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10314__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09107__C _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net318 _04003_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11970_ _05806_ _05814_ _05830_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__or3_1
X_10921_ net1461 net254 net487 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ net2209 net262 net491 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
X_13640_ clknet_leaf_92_clk net1277 net997 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13571_ clknet_leaf_61_clk top.a1.nextHex\[2\] net1110 vssd1 vssd1 vccd1 vccd1 _01379_
+ sky130_fd_sc_hd__dfrtp_1
X_10783_ net141 net2139 net372 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_51_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12522_ clknet_leaf_111_clk _00068_ net947 vssd1 vssd1 vccd1 vccd1 top.ramstore\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[16\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11404_ _05234_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__xnor2_4
X_12384_ _06157_ _06158_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11335_ top.a1.row1\[12\] _05127_ _05152_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11266_ top.lcd.nextState\[1\] _01382_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or2_1
XANTENNA__08177__A2 top.pc\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ net146 net1884 net441 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
X_13005_ clknet_leaf_112_clk _00551_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10224__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _01380_ _01427_ _01420_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08202__B _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__A1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07385__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net146 net2082 net445 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ net147 net2110 net446 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
XANTENNA__07137__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07105__Y _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ clknet_leaf_42_clk _01361_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12448__Q top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ clknet_leaf_73_clk _01294_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06310_ top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _01449_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08101__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07290_ _02393_ _02394_ _02403_ _02406_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nor4_2
XFILLER_0_127_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ wb.curr_state\[0\] _01407_ top.Wen wb.curr_state\[2\] _01400_ vssd1 vssd1
+ vccd1 vccd1 _00016_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_44_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06663__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06172_ top.a1.dataIn\[25\] vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold303 top.DUT.register\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 top.DUT.register\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 top.DUT.register\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 top.DUT.register\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 top.DUT.register\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold358 top.DUT.register\[13\]\[10\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 top.DUT.register\[12\]\[7\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _04915_ _04917_ _04914_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_4_3__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 _01553_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
Xfanout816 _04191_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_4_7__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout827 _01593_ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
X_09862_ _04494_ net360 net328 top.a1.dataIn\[20\] net363 vssd1 vssd1 vccd1 vccd1
+ _04856_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_2
Xfanout849 _05056_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_4
XANTENNA__07376__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ _03869_ _03906_ net317 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
Xhold1003 top.DUT.register\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ top.a1.dataIn\[13\] _04766_ _04792_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_
+ sky130_fd_sc_hd__a211o_1
Xhold1014 top.DUT.register\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 top.DUT.register\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1036 top.DUT.register\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 top.DUT.register\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _03082_ _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__xnor2_1
Xhold1058 top.DUT.register\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 top.a1.row2\[8\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07679__A1 _02795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _03734_ _03775_ _02716_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout453_A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07015__Y _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ net346 _02740_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ top.DUT.register\[11\]\[9\] net701 net558 top.DUT.register\[8\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout620_A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout718_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06508_ _01487_ _01489_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nor2_1
X_07488_ top.DUT.register\[26\]\[7\] net681 net669 top.DUT.register\[31\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06654__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09227_ net137 _04270_ _04275_ net133 _04274_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06439_ net810 _01527_ net808 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__and3_1
XANTENNA__10309__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09158_ _01778_ _02428_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _03219_ _03221_ _03223_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06406__A2 top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _03413_ _03449_ net286 net272 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ net65 net885 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_92_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08303__A _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 top.DUT.register\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 top.DUT.register\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net28 net862 net834 net1221 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__o22a_1
Xhold892 top.DUT.register\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10044__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net176 net2329 net451 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__mux2_1
XANTENNA__10979__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07119__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11953_ _05796_ _05797_ _05776_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08867__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10904_ net1846 net185 net407 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11884_ _05704_ _05739_ _05744_ _05735_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_67_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13623_ clknet_leaf_88_clk net1264 net1017 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06893__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10835_ net1446 net195 net494 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__mux2_1
XANTENNA__09788__B _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13554_ clknet_leaf_106_clk _01100_ net982 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10766_ net208 top.DUT.register\[25\]\[14\] net370 vssd1 vssd1 vccd1 vccd1 _00904_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ clknet_leaf_92_clk _00051_ net996 vssd1 vssd1 vccd1 vccd1 top.ramstore\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06645__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ clknet_leaf_114_clk _01031_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ net1459 net220 net498 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12436_ clknet_leaf_78_clk top.ru.next_FetchedData\[31\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11839__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12367_ _06146_ _06147_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output82_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ net900 _05127_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor2_1
XANTENNA__09309__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12298_ _06105_ net1118 _06104_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__and3b_1
X_11249_ _05124_ net1273 net402 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07358__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10889__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06790_ top.DUT.register\[29\]\[30\] net787 net718 top.DUT.register\[9\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08460_ net308 net302 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__or2_2
XFILLER_0_187_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07530__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07411_ top.a1.instruction\[26\] net854 _02527_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08391_ net287 _03376_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__nor2_1
XANTENNA__06884__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07342_ top.DUT.register\[15\]\[6\] net807 net803 top.DUT.register\[31\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08086__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ top.DUT.register\[23\]\[2\] net733 net761 top.DUT.register\[30\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a22o_1
XANTENNA__10129__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _02660_ net620 net1325 net887 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06224_ net1260 net1479 top.busy_o vssd1 vssd1 vccd1 vccd1 top.ru.next_dready sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold111 top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold144 top.ramaddr\[27\] vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 top.ramaddr\[28\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 top.ramaddr\[17\] vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 top.ramaddr\[15\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold199 top.DUT.register\[31\]\[10\] vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ net820 _04567_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__o21bai_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_8
Xfanout613 _06069_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 net626 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_4
XANTENNA__07349__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_4
Xfanout646 _01698_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08010__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _03820_ net454 net533 _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o211a_2
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10799__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _01684_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08410__X _03522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _01675_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
XANTENNA_fanout668_A _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ net818 _04336_ net816 top.pc\[11\] vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a2bb2o_1
X_06988_ top.DUT.register\[8\]\[20\] net593 net708 top.DUT.register\[7\]\[20\] _02104_
+ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08727_ _03788_ _03824_ net317 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13546__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ net1327 net859 net837 _03759_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07521__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09934__B1_N _04920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07609_ top.DUT.register\[22\]\[11\] net553 net636 top.DUT.register\[25\]\[11\] _02725_
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_194_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06875__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ net467 _03693_ _03688_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10620_ net240 net2158 net375 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XANTENNA__09401__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ net145 net1744 net428 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__mux2_1
XANTENNA__10039__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09026__B1 _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ net154 net2195 net505 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
X_13270_ clknet_leaf_105_clk _00816_ net982 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ net1320 net868 net832 _05942_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07588__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12152_ _06004_ _06011_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07052__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ net1232 net882 net848 top.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 _01182_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12083_ _05940_ _05941_ _05934_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a21o_1
XANTENNA__08810__A1_N net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ net1191 _05045_ net480 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10502__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12985_ clknet_leaf_58_clk _00531_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09501__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11936_ _05760_ _05751_ _05757_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__mux2_4
XFILLER_0_169_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07512__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11867_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13606_ clknet_leaf_74_clk _01147_ net1088 vssd1 vssd1 vccd1 vccd1 top.ramload\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818_ net1472 net240 net494 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
XANTENNA__09265__B1 _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ _05626_ net129 vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13537_ clknet_leaf_45_clk _01083_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10749_ net144 top.DUT.register\[24\]\[30\] net417 vssd1 vssd1 vccd1 vccd1 _00888_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09017__B1 _03102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13468_ clknet_leaf_17_clk _01014_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12419_ clknet_leaf_53_clk top.ru.next_FetchedData\[14\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13399_ clknet_leaf_112_clk _00945_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07579__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08240__A1 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__Q top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _03070_ _03072_ _03074_ _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_4_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11127__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06911_ _01943_ _02027_ net294 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__mux2_2
X_07891_ net353 _03004_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09630_ top.a1.instruction\[30\] net842 _04343_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10412__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06842_ top.DUT.register\[23\]\[27\] net730 net766 top.DUT.register\[11\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07751__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ top.DUT.register\[16\]\[29\] net723 net748 top.DUT.register\[1\]\[29\] _01889_
+ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a221o_1
X_09561_ net840 _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nor2_4
X_08512_ net469 _03608_ _03618_ net394 _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a221o_1
X_09492_ net840 _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__nor2_2
XFILLER_0_203_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07503__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09502__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _03428_ _03431_ net295 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06857__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06845__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08374_ _02562_ net458 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07325_ top.DUT.register\[5\]\[7\] net602 net778 top.DUT.register\[18\]\[7\] _02441_
+ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1060_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07256_ top.DUT.register\[7\]\[3\] net709 net749 top.DUT.register\[1\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XANTENNA__07282__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06207_ top.a1.halfData\[5\] _01426_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__nor2_2
XANTENNA__11479__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ _02289_ _02298_ _02301_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nor4_1
XFILLER_0_131_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout785_A _01534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout410 _04998_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
Xfanout421 _04994_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_6
XANTENNA_input9_X net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout443 net445 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_8
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_2
XANTENNA__09731__A1 _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout487 _05002_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_6
XANTENNA__10322__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ top.pc\[17\] _04445_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout498 net500 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_6
XANTENNA__07742__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ net813 _01626_ _04177_ _01620_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_87_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12770_ clknet_leaf_15_clk _00316_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11721_ _05543_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06848__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11652_ _05481_ _05489_ _05496_ _05498_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_37_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ net199 net2257 net422 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__A1 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ _05432_ _05433_ _05408_ _05410_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a211o_1
X_13322_ clknet_leaf_2_clk _00868_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire844 _01457_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_2
X_10534_ net213 top.DUT.register\[18\]\[13\] net426 vssd1 vssd1 vccd1 vccd1 _00679_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07273__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13253_ clknet_leaf_43_clk _00799_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ net227 net2027 net505 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__mux2_1
XANTENNA__11357__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12204_ top.a1.dataIn\[1\] _06063_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__xor2_1
XANTENNA__07025__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ clknet_leaf_106_clk _00730_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ net1418 net233 net515 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12135_ _05990_ _05992_ _05984_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07981__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _05901_ _05924_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a21bo_1
X_11017_ top.a1.data\[1\] net797 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__or2_1
XANTENNA__10232__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12968_ clknet_leaf_26_clk _00514_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _05735_ _05778_ _05779_ _05731_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a22oi_2
XANTENNA__06839__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ clknet_leaf_34_clk _00445_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13145__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12456__Q top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08880__B _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ top.DUT.register\[14\]\[14\] net792 net775 top.DUT.register\[2\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
X_08090_ _02174_ _03203_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__and2_1
XANTENNA__07264__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06681__A _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06472__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07041_ top.DUT.register\[16\]\[17\] net725 net761 top.DUT.register\[30\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a22o_1
Xclkload31 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_6
Xclkload42 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_8
XANTENNA__10407__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload53 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_6
Xclkload64 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_8
Xclkload75 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__clkinv_8
Xclkload86 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload97 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_2_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07783__Y _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ _04066_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__and3_2
XANTENNA__07972__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ _02958_ _02982_ _03009_ _03059_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_145_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10142__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ top.DUT.register\[21\]\[27\] net568 net544 top.DUT.register\[24\]\[27\] _02990_
+ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a221o_1
X_09613_ top.pc\[29\] _04614_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_207_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06825_ net324 _01941_ _01921_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__o21a_1
XFILLER_0_211_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09544_ net137 _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06756_ top.DUT.register\[15\]\[28\] net807 net589 top.DUT.register\[20\]\[28\] _01867_
+ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ _04497_ _04499_ _04495_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__o21ai_2
X_06687_ top.a1.instruction\[11\] _01486_ _01634_ top.a1.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 _01804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout533_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _03483_ _03536_ net313 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ net294 _02027_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout700_A _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12512__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07308_ top.DUT.register\[13\]\[1\] net791 net774 top.DUT.register\[2\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07255__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08452__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ net319 _03402_ _03400_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_210_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06463__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10317__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ _02349_ _02351_ _02353_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10250_ net147 net1366 net382 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__mux2_1
XANTENNA__07007__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ net1971 net145 net528 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout240 _04742_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
Xfanout273 _01858_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10052__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 _01800_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06518__B2 top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ net1131 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_198_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12822_ clknet_leaf_105_clk _00368_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13168__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ clknet_leaf_9_clk _00299_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11704_ _05534_ _05541_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ clknet_leaf_2_clk _00230_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11635_ _05492_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07246__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11566_ _05375_ _05399_ net248 vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ clknet_leaf_59_clk _00851_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06454__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ net147 net1801 net378 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__mux2_1
XANTENNA__10227__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11497_ _05321_ _05331_ _05356_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08205__B _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13236_ clknet_leaf_108_clk _00782_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10448_ net1405 net160 net511 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13167_ clknet_leaf_22_clk _00713_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ net1368 net168 net433 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07954__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _05949_ _05961_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__or2_1
XANTENNA__09317__A _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ clknet_leaf_118_clk _00644_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ _05892_ _05894_ _05884_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_127_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10897__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06610_ _01596_ _01726_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__nand2_2
X_07590_ top.DUT.register\[2\]\[15\] net685 net633 top.DUT.register\[27\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ top.a1.instruction\[22\] top.a1.instruction\[23\] net799 vssd1 vssd1 vccd1
+ vccd1 _01658_ sky130_fd_sc_hd__and3b_2
XFILLER_0_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08131__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06472_ top.DUT.register\[28\]\[0\] net739 net589 top.DUT.register\[20\]\[0\] _01571_
+ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a221o_1
X_09260_ top.pc\[9\] _02748_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__and2b_1
XANTENNA__07485__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08211_ net324 _02024_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__nor2_1
X_09191_ _01411_ _01753_ _04229_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__o21a_1
XANTENNA__06693__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ _03159_ _03208_ _03256_ _03258_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or4_1
XANTENNA__07237__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08073_ top.DUT.register\[22\]\[17\] net553 net648 top.DUT.register\[12\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a22o_1
XANTENNA__10137__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__B _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ top.DUT.register\[30\]\[18\] net760 net711 top.DUT.register\[25\]\[18\] _02140_
+ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09926__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1023_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _04040_ _04060_ net539 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21ai_1
Xhold15 top.a1.dataInTemp\[10\] vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 net110 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold37 top.a1.dataInTemp\[2\] vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ top.DUT.register\[5\]\[25\] net542 net630 top.DUT.register\[29\]\[25\] _03042_
+ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a221o_1
Xhold48 top.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 net74 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07857_ top.DUT.register\[15\]\[26\] net690 net542 top.DUT.register\[5\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout650_A _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__A0 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10600__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ top.DUT.register\[12\]\[31\] net736 net602 top.DUT.register\[5\]\[31\] _01924_
+ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07788_ _02903_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_203_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ _02024_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06739_ _01833_ _01854_ net826 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__mux2_4
XANTENNA_fanout915_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09897__A _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ net841 _02589_ net618 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09870__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ net462 _03497_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06592__Y _01709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _04412_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11420_ top.a1.dataIn\[27\] _05251_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__xor2_1
XANTENNA__12221__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_X clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _05206_ _05213_ _05214_ net843 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__or4b_1
XFILLER_0_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ net2266 net208 net521 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ _05147_ _05150_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_111_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13021_ clknet_leaf_119_clk _00567_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09925__A1 _03977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ net218 net1850 net382 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XANTENNA__07936__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ top.DUT.register\[7\]\[13\] net214 net525 vssd1 vssd1 vccd1 vccd1 _00327_
+ sky130_fd_sc_hd__mux2_1
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09137__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
Xfanout1024 net1030 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1035 net1038 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
X_10095_ net219 net2264 net387 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
Xfanout1068 net1072 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1121 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_4
XFILLER_0_89_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08900__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ clknet_leaf_60_clk _01377_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10510__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ clknet_leaf_39_clk _00351_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ clknet_leaf_65_clk _01310_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10997_ net1169 _05017_ net480 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12736_ clknet_leaf_14_clk _00282_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07467__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06675__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ clknet_leaf_5_clk _00213_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07219__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ _05442_ net207 _05474_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__o22ai_4
XANTENNA__12212__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12598_ clknet_leaf_105_clk _00144_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08967__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11549_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold507 top.pad.keyCode\[2\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 top.DUT.register\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 top.DUT.register\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08650__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13219_ clknet_leaf_35_clk _00765_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11577__A top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07927__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _03806_ _03856_ _03154_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a21o_1
X_07711_ _02448_ _02611_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nand2b_1
XANTENNA_wire337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ _03703_ _03790_ net295 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08352__B1 _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07642_ top.DUT.register\[18\]\[8\] net661 net637 top.DUT.register\[25\]\[8\] _02758_
+ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a221o_1
XANTENNA__09954__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ _02346_ _02688_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08104__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09312_ top.pc\[12\] _04344_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or2_1
X_06524_ top.a1.instruction\[29\] _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__and2_1
XANTENNA__08655__A1 _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07458__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__B2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09510__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06666__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ net137 _04284_ _04290_ net822 vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o22a_1
X_06455_ top.DUT.register\[29\]\[0\] net785 net585 top.DUT.register\[24\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout231_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06386_ top.pad.button_control.r_counter\[5\] top.pad.button_control.r_counter\[6\]
+ top.pad.button_control.r_counter\[7\] vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o21a_1
X_09174_ _01411_ _01753_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08125_ top.DUT.register\[3\]\[16\] net691 net683 top.DUT.register\[2\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07091__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ top.DUT.register\[23\]\[23\] net565 net672 top.DUT.register\[19\]\[23\] _03172_
+ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_186_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout698_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ top.DUT.register\[8\]\[19\] net592 net584 top.DUT.register\[24\]\[19\] _02123_
+ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a221o_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__07918__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08591__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ _02905_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_90_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ top.DUT.register\[25\]\[24\] net638 net625 top.DUT.register\[16\]\[24\] _03025_
+ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a221o_1
X_08889_ net904 top.pc\[26\] _03978_ _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net1367 net265 net487 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__mux2_1
XANTENNA__10330__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ net1424 net241 net490 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ clknet_leaf_61_clk top.a1.nextHex\[1\] net1110 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10782_ net143 net2071 net373 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ clknet_leaf_92_clk _00067_ net996 vssd1 vssd1 vccd1 vccd1 top.ramstore\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06657__B1 _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12452_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[15\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08036__A _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _05236_ _05246_ net478 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__and3_2
X_12383_ net1278 _06155_ net815 vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11334_ net1202 net843 _05201_ net1115 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ net901 top.lcd.nextState\[1\] top.lcd.nextState\[0\] _05130_ vssd1 vssd1
+ vccd1 vccd1 _05136_ sky130_fd_sc_hd__and4_1
XANTENNA__10505__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__Y _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ clknet_leaf_3_clk _00550_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10216_ net147 top.DUT.register\[8\]\[29\] net438 vssd1 vssd1 vccd1 vccd1 _00375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ _01420_ _05096_ _05101_ _05100_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a31o_1
XANTENNA__11181__A2 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ net149 net2173 net442 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA__08819__B1_N _03229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10078_ net151 net2135 net448 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
XANTENNA__10240__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ clknet_leaf_42_clk _01360_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13768_ clknet_leaf_66_clk _01293_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__B2 _03739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09330__A top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ clknet_leaf_22_clk _00265_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07769__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ clknet_leaf_62_clk _01232_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06240_ wb.curr_state\[0\] top.Ren _01408_ wb.curr_state\[1\] net925 vssd1 vssd1
+ vccd1 vccd1 _00015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_170_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13664__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06171_ top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 top.DUT.register\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07785__A _01920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold315 top.DUT.register\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 top.DUT.register\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 top.DUT.register\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold348 top.DUT.register\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ top.pc\[27\] _04606_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__nor2_1
Xhold359 top.DUT.register\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10415__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 _01553_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
X_09861_ _04853_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout817 _04191_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
Xfanout839 _03295_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_0_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08812_ _03328_ _03331_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_181_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1004 top.DUT.register\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ net818 _04370_ _04790_ _04791_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__o22ai_1
Xhold1015 top.DUT.register\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 top.DUT.register\[27\]\[6\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _03157_ _03822_ _03155_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09505__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1037 top.DUT.register\[16\]\[6\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 top.DUT.register\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 top.DUT.register\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout181_A _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _02640_ _02717_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _02305_ _02740_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_200_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08628__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ top.DUT.register\[1\]\[9\] net705 net574 top.DUT.register\[7\]\[9\] _02672_
+ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_196_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08628__B2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06639__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ _01487_ _01491_ _01610_ _01617_ _01623_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__o311a_1
X_07487_ top.DUT.register\[8\]\[7\] net558 net641 top.DUT.register\[9\]\[7\] _02603_
+ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_46_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09226_ top.pc\[6\] _04254_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06438_ net811 _01518_ _01536_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__and3_1
XANTENNA__07851__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09157_ net367 _01643_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__nor2_1
XANTENNA__13334__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06369_ top.d_ready _01487_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07064__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ top.DUT.register\[23\]\[22\] net565 net648 top.DUT.register\[12\]\[22\] _03224_
+ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a221o_1
XANTENNA__08290__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ _03485_ _03538_ _03564_ net272 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06811__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ _02131_ _03152_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_92_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10325__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 top.DUT.register\[23\]\[29\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold871 top.DUT.register\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 top.DUT.register\[14\]\[5\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net27 net851 net850 net1902 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a22o_1
Xhold893 top.DUT.register\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net181 net1791 net451 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06590__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10060__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _05768_ _05799_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06477__C top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10903_ net2230 net189 net406 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
X_11883_ top.a1.dataIn\[5\] _05740_ _05741_ _05742_ vssd1 vssd1 vccd1 vccd1 _05744_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_196_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13622_ clknet_leaf_75_clk net1160 net1083 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
X_10834_ net2242 net199 net493 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ clknet_leaf_7_clk _01099_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ net213 net2192 net370 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08095__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12504_ clknet_leaf_78_clk net34 net1080 vssd1 vssd1 vccd1 vccd1 top.testpc.en_latched
+ sky130_fd_sc_hd__dfrtp_2
X_13484_ clknet_leaf_3_clk _01030_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07842__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10696_ net1654 net227 net497 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ clknet_leaf_74_clk top.ru.next_FetchedData\[30\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[30\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12366_ _01404_ _06145_ net814 vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ top.lcd.nextState\[3\] net900 _05127_ top.lcd.nextState\[4\] vssd1 vssd1
+ vccd1 vccd1 _05185_ sky130_fd_sc_hd__or4b_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10235__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ top.lcd.cnt_20ms\[16\] top.lcd.cnt_20ms\[15\] _06101_ vssd1 vssd1 vccd1 vccd1
+ _06105_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_73_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ net871 _05111_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ net138 _04721_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12459__Q top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07410_ _01630_ _01803_ _02526_ net400 net857 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a221o_1
X_08390_ net283 _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__and2_1
XANTENNA__09807__B1 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09060__A _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07341_ _02451_ _02453_ _02455_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__or4_2
XANTENNA__08086__A2 _03202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07294__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ _02376_ _02385_ _02386_ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__nor4_2
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ _02819_ net620 net1184 net888 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09015__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06223_ top.busy_o top.ru.state\[4\] vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__and2b_1
XANTENNA__07786__Y _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07046__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _01354_ vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold123 top.a1.row1\[122\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 top.a1.row1\[17\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 top.pad.button_control.noisy vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10145__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 top.ramaddr\[6\] vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold167 top.ramaddr\[8\] vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold178 top.ramstore\[20\] vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _04576_ net360 net329 top.a1.dataIn\[25\] net364 vssd1 vssd1 vccd1 vccd1
+ _04902_ sky130_fd_sc_hd__a221o_1
Xhold189 top.ramstore\[24\] vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout603 _01538_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_4
XFILLER_0_186_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout614 _04728_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11765__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _01701_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_4
Xfanout647 _01696_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
X_09844_ _04192_ _04838_ _04839_ _04835_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout658 _01691_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
XANTENNA__08010__A2 _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _01684_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_8
X_09775_ net223 top.DUT.register\[1\]\[10\] net390 vssd1 vssd1 vccd1 vccd1 _00132_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout563_A _01673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ top.DUT.register\[14\]\[20\] net793 net720 top.DUT.register\[26\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08726_ _03334_ _03338_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08657_ net902 top.pc\[15\] net537 _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout730_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07608_ top.DUT.register\[28\]\[11\] net656 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_194_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _03691_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__nand2_1
XANTENNA__06594__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07539_ top.DUT.register\[11\]\[13\] net699 net544 top.DUT.register\[24\]\[13\] _02655_
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08077__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11081__A1 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10__f_clk_X clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ net147 net1858 net426 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__mux2_1
XANTENNA__07285__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _04244_ _04246_ _04257_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10481_ net159 net1940 net505 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09026__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ net1274 net867 net832 _05964_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _06004_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10055__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ net1276 net878 net846 top.ramstore\[20\] vssd1 vssd1 vccd1 vccd1 _01181_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12082_ _05940_ _05941_ _05929_ _05930_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__o2bb2a_1
Xhold690 top.DUT.register\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
X_11033_ net864 _05043_ _05044_ net869 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1
+ _05045_ sky130_fd_sc_hd__a32o_1
XANTENNA__08001__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A _02519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ clknet_leaf_33_clk _00530_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ _05785_ _05786_ _05794_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a21o_2
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09799__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11866_ _05693_ _05725_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13605_ clknet_leaf_74_clk _01146_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramload\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_205_Right_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ _04183_ net616 _04973_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_31_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09265__A1 _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08068__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ _01399_ _05654_ _05655_ _05656_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_31_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13536_ clknet_leaf_12_clk _01082_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07276__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ net147 net2286 net414 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13467_ clknet_leaf_5_clk _01013_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09017__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ net161 net2228 net420 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07028__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12418_ clknet_leaf_53_clk top.ru.next_FetchedData\[13\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[13\] sky130_fd_sc_hd__dfrtp_4
X_13398_ clknet_leaf_105_clk _00944_ net981 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12349_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[1\]
+ top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a21o_1
XANTENNA__09039__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06910_ _01984_ _02026_ net319 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07890_ net353 _03004_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__nand2_1
XANTENNA__07200__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06841_ top.DUT.register\[16\]\[27\] net723 net596 top.DUT.register\[6\]\[27\] _01957_
+ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ top.a1.instruction\[26\] net842 net618 vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a21oi_1
X_06772_ top.DUT.register\[14\]\[29\] net792 net734 top.DUT.register\[12\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ _02695_ net458 _03615_ net474 _03609_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a221o_1
X_09491_ net841 _01777_ net618 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08442_ _03427_ _03435_ net287 vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ net476 _02560_ _02561_ net396 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07267__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ top.DUT.register\[12\]\[7\] net737 net729 top.DUT.register\[10\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a22o_1
XANTENNA__11063__A1 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07806__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07255_ top.DUT.register\[15\]\[3\] net806 net802 top.DUT.register\[31\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout311_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1053_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A _05001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06206_ _01423_ _01424_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__and2_1
XANTENNA__07019__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07186_ top.DUT.register\[22\]\[11\] net605 net720 top.DUT.register\[26\]\[11\] _02302_
+ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a221o_1
XANTENNA__08231__A2 _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _01629_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
Xfanout411 _04998_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06793__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net425 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _04984_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_6
Xfanout455 _04737_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
Xfanout477 _01729_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
X_09827_ top.pc\[16\] _04425_ _04817_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_129_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09731__A2 _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout488 _05002_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout945_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_8
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__inv_2
XANTENNA__06876__X _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13767__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08709_ _03806_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09689_ net907 _01480_ _04708_ net1102 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ _05547_ _05548_ _05579_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13865__1126 vssd1 vssd1 vccd1 vccd1 _13865__1126/HI net1126 sky130_fd_sc_hd__conb_1
X_11651_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07258__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__A1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net205 net1549 net424 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__A2 _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11582_ _05438_ _05439_ _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ clknet_leaf_28_clk _00867_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10533_ net216 net1515 net426 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9__f_clk_X clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_30_clk _00798_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10464_ net228 net2201 net507 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12203_ top.a1.dataIn\[1\] _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_114_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13183_ clknet_leaf_22_clk _00729_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ net1554 net238 net516 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
X_12134_ _05987_ _05989_ _05990_ _05992_ _05984_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__o2111a_1
XANTENNA__06784__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10513__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ _05879_ _05899_ _05900_ _05876_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__o2bb2a_1
X_11016_ top.a1.dataInTemp\[5\] net798 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07107__B _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12967_ clknet_leaf_49_clk _00513_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net125 _05759_ _05769_ _05734_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a211o_1
XFILLER_0_197_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08219__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ clknet_leaf_11_clk _00444_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11849_ _05682_ _05686_ _05668_ _05672_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ clknet_leaf_20_clk _01065_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_8
Xclkload21 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_6
X_07040_ top.DUT.register\[10\]\[17\] net727 net749 top.DUT.register\[1\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload32 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload43 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload43/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__inv_16
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload65 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__bufinv_16
Xclkload76 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload87 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_16
Xclkload98 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_2_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08991_ net465 _04068_ _04075_ _02879_ _04073_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__o221a_1
XANTENNA__06775__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ _03032_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or2_1
XANTENNA__10423__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12204__A top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ top.DUT.register\[19\]\[27\] net671 net643 top.DUT.register\[10\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09612_ top.pc\[29\] _04614_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__and2_1
X_06824_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_178_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09543_ _04571_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__xnor2_1
X_06755_ top.DUT.register\[27\]\[28\] net771 net716 top.DUT.register\[9\]\[28\] _01866_
+ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout261_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07488__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _04506_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09232__B _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06686_ top.a1.instruction\[17\] net824 _01640_ top.a1.instruction\[25\] vssd1 vssd1
+ vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ net321 _02468_ _02490_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_82_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout526_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ net294 _02112_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08988__A0 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinvlp_4
X_07307_ top.DUT.register\[28\]\[1\] net740 net583 top.DUT.register\[4\]\[1\] _02423_
+ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08287_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__inv_2
XANTENNA__06226__C_N net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07660__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ top.DUT.register\[26\]\[8\] net721 net586 top.DUT.register\[24\]\[8\] _02354_
+ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07169_ _02245_ _02285_ net315 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
X_10180_ net2318 net148 net525 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 _04742_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_1
XANTENNA__09165__B1 _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 _04756_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_199_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout274 net276 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
Xfanout285 _01800_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
Xfanout296 _01774_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
X_13870_ net1130 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_198_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07191__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ clknet_leaf_100_clk _00367_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07479__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ clknet_leaf_114_clk _00298_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11703_ _05532_ _05550_ _05531_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12683_ clknet_leaf_4_clk _00229_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12224__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ _05493_ _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10508__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ _05421_ _05422_ _05397_ _05420_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_25_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ clknet_leaf_37_clk _00850_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07651__A0 _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12487__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10516_ net153 net2040 net379 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__mux2_1
X_11496_ _05302_ _05317_ _05353_ _05330_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__or4b_1
X_13235_ clknet_leaf_111_clk _00781_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net1397 net162 net512 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08061__X _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ clknet_leaf_95_clk _00712_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net1573 net173 net430 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
X_12117_ _05967_ _05968_ _05971_ _05973_ _05976_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10243__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ clknet_leaf_27_clk _00643_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__B _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ _05871_ _05903_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08648__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07182__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__X _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _01646_ _01649_ _01656_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__and3_4
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12467__Q top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06471_ top.DUT.register\[23\]\[0\] net731 _01585_ _01587_ vssd1 vssd1 vccd1 vccd1
+ _01588_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08210_ net278 _03317_ _03325_ net270 _03310_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07788__A _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__B2 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ _04239_ _04240_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06692__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _03183_ _03232_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or2_1
XANTENNA__10418__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08072_ top.DUT.register\[24\]\[17\] net545 _03188_ vssd1 vssd1 vccd1 vccd1 _03189_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07642__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06996__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ top.DUT.register\[10\]\[18\] net726 net725 top.DUT.register\[16\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06748__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10153__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864__1125 vssd1 vssd1 vccd1 vccd1 _13864__1125/HI net1125 sky130_fd_sc_hd__conb_1
X_08974_ _04040_ _04060_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1016_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 top.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 top.a1.data\[6\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ top.DUT.register\[22\]\[25\] net555 net638 top.DUT.register\[25\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a22o_1
Xhold38 top.a1.dataInTemp\[3\] vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold49 top.ramstore\[26\] vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ top.DUT.register\[6\]\[26\] net577 net624 top.DUT.register\[16\]\[26\] _02972_
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a221o_1
XFILLER_0_194_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08370__A1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ top.DUT.register\[21\]\[31\] net610 net607 top.DUT.register\[22\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
X_07787_ _01919_ _02901_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06920__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ net840 _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_27_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06738_ _01834_ _01853_ net826 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _04488_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06669_ top.DUT.register\[21\]\[1\] net570 net633 top.DUT.register\[27\]\[1\] _01785_
+ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ net464 _03519_ _03517_ _03512_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07881__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _04408_ _04413_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_81_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08339_ _02845_ _03418_ _02842_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08425__A2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__A1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07985__X _03102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ top.a1.row1\[15\] _05152_ _05184_ net900 _05210_ vssd1 vssd1 vccd1 vccd1
+ _05214_ sky130_fd_sc_hd__a221o_1
XANTENNA__07633__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ top.DUT.register\[11\]\[13\] net212 net521 vssd1 vssd1 vccd1 vccd1 _00455_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06987__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ _05147_ _05150_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_111_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13020_ clknet_leaf_18_clk _00566_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ net219 net1949 net383 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XANTENNA__09925__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10063__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1003 net1021 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_4
X_10163_ net2123 net218 net525 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XANTENNA__07209__Y _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 net1020 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_2
Xfanout1025 net1030 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_206_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1036 net1038 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_2
XANTENNA_input37_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1050 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_2
X_10094_ net226 net1876 net386 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
Xfanout1058 net1073 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_2
Xfanout1069 net1072 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07164__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13853_ clknet_leaf_60_clk _01376_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08900__A3 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ clknet_leaf_30_clk _00350_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10996_ top.a1.dataIn\[0\] net870 _05014_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_
+ sky130_fd_sc_hd__a22o_1
X_13784_ clknet_leaf_65_clk _01309_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12735_ clknet_leaf_23_clk _00281_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07872__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ clknet_leaf_15_clk _00212_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07401__A _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11617_ _05438_ _05439_ _05442_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__and3_1
XANTENNA__10238__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ clknet_leaf_100_clk _00143_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11548_ _05383_ _05405_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06978__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 top.DUT.register\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 top.DUT.register\[16\]\[5\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ top.a1.dataIn\[17\] _05305_ _05330_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ clknet_leaf_12_clk _00764_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13149_ clknet_leaf_119_clk _00695_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1208 top.ramstore\[22\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
X_07710_ _02745_ _02773_ _02825_ _02826_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__or4_1
X_08690_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__inv_2
XANTENNA__10701__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__B2 _03465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ top.DUT.register\[15\]\[8\] net689 net657 top.DUT.register\[28\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
XANTENNA__06902__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07572_ net829 net331 _02669_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_66_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09311_ top.pc\[12\] _04344_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__and2_1
XANTENNA__09350__X _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06523_ _01486_ _01634_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_157_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ _04285_ _04288_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ top.DUT.register\[21\]\[0\] net609 net735 top.DUT.register\[12\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13008__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09173_ _01410_ net853 _04225_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06385_ top.pad.button_control.r_counter\[10\] top.pad.button_control.r_counter\[9\]
+ top.pad.button_control.r_counter\[7\] top.pad.button_control.r_counter\[5\] vssd1
+ vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__nand4_1
XANTENNA__10148__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ _03234_ _03236_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__or3_1
XANTENNA__09937__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07615__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06969__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ top.DUT.register\[1\]\[23\] net704 net695 top.DUT.register\[30\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_186_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ top.DUT.register\[9\]\[19\] net715 net758 top.DUT.register\[2\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
XANTENNA__09238__A _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A _01551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08591__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08591__B2 _03695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _02931_ _04024_ _02929_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_90_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10611__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ top.DUT.register\[31\]\[24\] net670 net661 top.DUT.register\[18\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a22o_1
X_08888_ _03955_ _03977_ net539 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o21a_1
X_07839_ _02954_ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ net614 _04982_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ _02068_ net840 _04524_ _04526_ _04527_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10781_ net149 net2225 net370 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06657__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12520_ clknet_leaf_76_clk _00066_ net1082 vssd1 vssd1 vccd1 vccd1 top.ramstore\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12451_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[14\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[14\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10058__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ top.a1.dataIn\[31\] _05231_ _05259_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07606__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ top.pad.button_control.r_counter\[14\] top.pad.button_control.r_counter\[13\]
+ _06153_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3_1
X_11333_ _05192_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ top.a1.row2\[0\] _05132_ _05134_ top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1
+ _05135_ sky130_fd_sc_hd__a22o_1
X_13003_ clknet_leaf_6_clk _00549_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ net152 net1760 net440 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XANTENNA__08031__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _01379_ net907 _01427_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__mux2_1
XANTENNA__08987__A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07385__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _04932_ net1537 net444 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
XANTENNA__06593__A0 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10521__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ net155 net2100 net446 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07137__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload2_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ clknet_leaf_42_clk _01359_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08098__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13767_ clknet_leaf_66_clk _01292_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_10979_ net1600 net148 net481 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__B2 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__Y _02519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ clknet_leaf_95_clk _00264_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09330__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07845__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13863__1124 vssd1 vssd1 vccd1 vccd1 _13863__1124/HI net1124 sky130_fd_sc_hd__conb_1
X_13698_ clknet_leaf_62_clk _01231_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ clknet_leaf_26_clk _00195_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06170_ top.a1.dataIn\[19\] vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold305 top.DUT.register\[4\]\[4\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 top.DUT.register\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold327 top.DUT.register\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 top.DUT.register\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 top.DUT.register\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout807 _01553_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08022__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _04843_ _04846_ _04852_ _04192_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a31o_1
Xfanout818 _04170_ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_2
Xfanout829 _01592_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_4
XANTENNA__08573__A1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ _03183_ net459 _03903_ net395 _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a221o_1
XANTENNA__09770__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _04378_ net362 _04769_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_181_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 top.DUT.register\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1016 top.DUT.register\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 top.pad.button_control.r_counter\[6\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ net1322 net859 net836 _03839_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a22o_1
Xhold1038 top.DUT.register\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__B _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10431__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1049 top.DUT.register\[23\]\[4\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A2 _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ _03764_ _03766_ _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_163_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout174_A _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07624_ _02305_ _02740_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_200_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ top.DUT.register\[22\]\[9\] net554 net649 top.DUT.register\[12\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09825__A1 _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_clk_X clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ top.a1.instruction\[14\] _01487_ _01610_ vssd1 vssd1 vccd1 vccd1 _01623_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07486_ top.DUT.register\[2\]\[7\] net686 net649 top.DUT.register\[12\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08137__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07300__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ _04261_ _04271_ _04272_ _04273_ net822 vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_101_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06437_ top.a1.instruction\[19\] net830 _01552_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__and3_4
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09156_ net400 _04171_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06368_ _01488_ _01490_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__nor2_1
X_08107_ top.DUT.register\[7\]\[22\] net573 net624 top.DUT.register\[16\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09087_ _03927_ _03945_ _03970_ _03987_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10606__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06299_ net1324 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[25\] sky130_fd_sc_hd__and2_1
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _02131_ _03152_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold850 top.pad.button_control.r_counter\[4\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 top.DUT.register\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 top.DUT.register\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 top.DUT.register\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 top.DUT.register\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07367__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ net186 net2202 net450 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__mux2_1
XANTENNA__08564__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__B2 _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__X _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ net230 net1885 net452 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__mux2_1
XANTENNA__10341__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _05768_ _05799_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_106_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09134__C top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ net2155 net191 net406 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
X_11882_ _05741_ _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13621_ clknet_leaf_75_clk net1289 net1084 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
X_10833_ net1513 net206 net495 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09150__B _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13552_ clknet_leaf_116_clk _01098_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10764_ net216 net1686 net370 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XANTENNA__07827__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12503_ clknet_leaf_76_clk _00050_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ clknet_leaf_6_clk _01029_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net1380 net229 net498 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12434_ clknet_leaf_78_clk top.ru.next_FetchedData\[29\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12365_ _01404_ _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10516__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_101_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11316_ net906 _05148_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__nor2_1
X_12296_ top.lcd.cnt_20ms\[15\] top.lcd.cnt_20ms\[14\] _06100_ top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__a31o_1
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11247_ _05123_ net1253 net403 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XANTENNA__08004__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _01332_ _01334_ _01468_ _01477_ _01335_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a311oi_1
XANTENNA__10251__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net222 net2011 net443 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08858__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07530__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13819_ clknet_leaf_71_clk _01344_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06684__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__B2 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ top.DUT.register\[6\]\[6\] net598 net594 top.DUT.register\[8\]\[6\] _02456_
+ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a221o_1
XANTENNA__07818__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ top.DUT.register\[12\]\[3\] net736 net768 top.DUT.register\[11\]\[3\] _02387_
+ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ _02739_ net620 net1194 net887 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__a2bb2o_1
X_06222_ _00008_ top.a1.nextHex\[7\] vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[4\] sky130_fd_sc_hd__or2_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10426__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold102 top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 top.a1.row1\[121\] vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold124 top.ramstore\[3\] vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 top.a1.row2\[25\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 top.a1.row1\[13\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top.DUT.register\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold179 top.ramaddr\[13\] vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09912_ _04897_ _04898_ _04899_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_74_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_4
XFILLER_0_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout615 _04728_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_2
XANTENNA__07349__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout626 _01705_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09743__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _04836_ _04837_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nor2_1
Xfanout637 _01701_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08420__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 _01696_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_4
XANTENNA_fanout291_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 net662 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA__10161__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ top.DUT.register\[3\]\[20\] net782 net600 top.DUT.register\[5\]\[20\] _02102_
+ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a221o_1
X_09774_ _03646_ net454 net533 _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o211a_2
XANTENNA__07036__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ _03158_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_198_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout556_A net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _03742_ _03746_ _03753_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or4b_4
XFILLER_0_178_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__A2 _02637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07470__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ top.DUT.register\[7\]\[11\] net573 net672 top.DUT.register\[19\]\[11\] _02723_
+ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ _02824_ _03690_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout723_A _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07538_ top.DUT.register\[1\]\[13\] net703 net556 top.DUT.register\[8\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a22o_1
XANTENNA__07809__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07469_ _02576_ _02585_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09208_ _04244_ _04246_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__o21a_1
X_10480_ net165 net2178 net508 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__RESET_B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__A0 _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ net913 _01595_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or2_4
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10336__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _06001_ _06005_ _06002_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06796__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ net1211 net879 net847 top.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 _01180_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _05940_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__nand2_1
Xhold680 top.DUT.register\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08537__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold691 top.DUT.register\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ top.a1.data\[5\] net796 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__or2_1
XANTENNA__08537__B2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862__1123 vssd1 vssd1 vccd1 vccd1 _13862__1123/HI net1123 sky130_fd_sc_hd__conb_1
XANTENNA__10071__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12983_ clknet_leaf_107_clk _00529_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11934_ _05785_ _05786_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07512__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11865_ _05693_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__and2b_1
XANTENNA__06720__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13839__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ clknet_leaf_55_clk _01145_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramload\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_184_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10816_ net142 net1780 net412 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11796_ _05655_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09265__A2 _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13535_ clknet_leaf_23_clk _01081_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ net150 net1927 net415 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ net162 net1749 net420 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XANTENNA__09017__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13466_ clknet_leaf_15_clk _01012_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12417_ clknet_leaf_53_clk top.ru.next_FetchedData\[12\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[12\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10246__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ clknet_leaf_100_clk _00943_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07579__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[2\]
+ top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__and3_1
XANTENNA__06787__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_206_Left_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12279_ net1182 _06091_ _06093_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_56_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11127__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__Y _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ top.DUT.register\[5\]\[27\] net600 net726 top.DUT.register\[10\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ top.DUT.register\[26\]\[29\] net719 net588 top.DUT.register\[20\]\[29\] _01887_
+ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a221o_1
X_08510_ _03355_ _03569_ _03607_ _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_160_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ _04519_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08700__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07503__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _02832_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ _01801_ _03484_ net289 vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_2
XFILLER_0_92_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06982__X _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ top.DUT.register\[25\]\[7\] net713 _02439_ vssd1 vssd1 vccd1 vccd1 _02440_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout137_A _04208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06205_ top.a1.halfData\[5\] _01424_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10156__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ top.DUT.register\[31\]\[11\] net800 net756 top.DUT.register\[3\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout304_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06778__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _01629_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_2
Xfanout412 _04998_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_6
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_8
Xfanout445 _04971_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_4
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__B1 top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 _04737_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_4
X_09826_ net202 net1750 net390 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__mux2_1
Xfanout467 _03363_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
Xfanout478 _05263_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_2
Xfanout489 net492 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07742__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net813 _01626_ _01619_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_198_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06969_ top.DUT.register\[13\]\[21\] net789 net725 top.DUT.register\[16\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ _03107_ _03805_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _04695_ _04702_ _04705_ _04707_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__or4_1
X_08639_ _02720_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11650_ _05508_ _05510_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ net210 net2342 net422 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11581_ _05402_ _05403_ _05434_ _05440_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a32o_1
XFILLER_0_193_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ net220 net1988 net427 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__mux2_1
XANTENNA__07500__Y _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13320_ clknet_leaf_25_clk _00866_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ clknet_leaf_35_clk _00797_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10066__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ net234 net1529 net507 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08758__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _06059_ _06060_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__a21o_1
XANTENNA__08758__B2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ clknet_leaf_40_clk _00728_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08612__X _03716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ net1441 net245 net515 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XANTENNA__06769__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__B1 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _05987_ _05989_ _05990_ _05992_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07981__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _05901_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__nand2_1
X_11015_ net1390 _05031_ net480 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
XANTENNA__07194__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 net992 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09014__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06941__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12966_ clknet_leaf_19_clk _00512_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _05758_ _05759_ _05769_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12897_ clknet_leaf_43_clk _00443_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08219__B _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11848_ _05674_ _05686_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nor2_1
XANTENNA__09029__A2_N _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ _05629_ _05630_ _05638_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ clknet_leaf_94_clk _01064_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload11 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__06472__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload22 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_8
X_13449_ clknet_leaf_27_clk _00995_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload33 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload44 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08749__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload55 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__inv_16
XANTENNA__09946__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload66 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload77 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload88 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__inv_6
Xclkload99 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload99/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10704__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ net287 net275 _02517_ _03459_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _03056_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__nand2_2
XFILLER_0_167_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07872_ top.DUT.register\[20\]\[27\] net560 net659 top.DUT.register\[18\]\[27\] _02988_
+ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a221o_1
XANTENNA__07185__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__A1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net136 _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nor2_1
X_06823_ _01930_ _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nor2_4
XFILLER_0_211_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_178_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09542_ _04550_ _04551_ _04552_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__o21ai_2
X_06754_ top.DUT.register\[4\]\[28\] net582 net757 top.DUT.register\[3\]\[28\] _01870_
+ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06685_ net286 _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__or2_1
X_09473_ _04488_ _04489_ _04490_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_90_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09784__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08424_ net303 _03534_ _03529_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _02562_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_82_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout421_A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07306_ top.DUT.register\[29\]\[1\] net787 net709 top.DUT.register\[7\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout519_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13861__1122 vssd1 vssd1 vccd1 vccd1 _13861__1122/HI net1122 sky130_fd_sc_hd__conb_1
Xclkload5 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_61_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ net296 net356 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08145__A _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07237_ top.DUT.register\[12\]\[8\] net736 net728 top.DUT.register\[10\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
XANTENNA__06463__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ net300 _02284_ _02265_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__A1 top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ top.DUT.register\[20\]\[15\] net590 net586 top.DUT.register\[24\]\[15\] _02215_
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a221o_1
Xfanout220 _04781_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_1
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 _04775_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout242 _04742_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12711__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 net256 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 _04744_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07176__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09737__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_1
XFILLER_0_199_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout286 _01775_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XFILLER_0_198_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout297 net300 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
X_09809_ top.pc\[15\] _04410_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2_1
XANTENNA__06923__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ clknet_leaf_99_clk _00366_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ clknet_leaf_20_clk _00297_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__C1 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10483__A0 _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11702_ _05558_ _05561_ _05556_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__o21bai_1
X_12682_ clknet_leaf_117_clk _00228_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11633_ _05454_ _05465_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__and4b_1
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10235__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06782__B _01898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11564_ _05422_ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__or2_1
XANTENNA__07100__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09640__A2 _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ clknet_leaf_109_clk _00849_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07651__A1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10515_ net156 net1779 net379 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__mux2_1
XANTENNA__06454__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11495_ _05327_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ net1399 net166 net512 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__mux2_1
X_13234_ clknet_leaf_107_clk _00780_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10524__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13165_ clknet_leaf_115_clk _00711_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10377_ net1975 net177 net431 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07954__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ _05971_ _05973_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__or3_1
X_13096_ clknet_leaf_24_clk _00642_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12452__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _05876_ _05901_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06914__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ clknet_leaf_101_clk _00495_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_72_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08131__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06470_ top.DUT.register\[31\]\[0\] net800 net749 top.DUT.register\[1\]\[0\] _01547_
+ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06973__A _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06693__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08140_ _03256_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload100 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload100/X sky130_fd_sc_hd__clkbuf_8
X_08071_ top.DUT.register\[11\]\[17\] net700 net640 top.DUT.register\[9\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a22o_1
X_07022_ top.DUT.register\[14\]\[18\] net792 net758 top.DUT.register\[2\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_157_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10434__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09395__B2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07945__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _04054_ _04055_ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 _01176_ vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 top.a1.data\[5\] vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _03034_ _03036_ _03038_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__or4_1
Xhold39 top.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09524__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ top.DUT.register\[14\]\[26\] net664 net652 top.DUT.register\[17\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout371_A _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ top.DUT.register\[30\]\[31\] net762 net582 top.DUT.register\[4\]\[31\] _01922_
+ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_166_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07786_ _01919_ _02901_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_84_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09525_ top.a1.instruction\[24\] net842 net618 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a21oi_1
X_06737_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__C1 _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout636_A _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ top.DUT.register\[7\]\[1\] net575 net551 top.DUT.register\[4\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a22o_1
X_09456_ _04489_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08407_ _02841_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ net350 _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__xnor2_1
X_06599_ top.a1.instruction\[22\] top.a1.instruction\[23\] _01714_ _01715_ vssd1 vssd1
+ vccd1 vccd1 _01716_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout803_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10217__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ net474 net277 _03451_ _03445_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a31o_1
XANTENNA__09083__B1 _03772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _02196_ _02245_ net315 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_175_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10300_ net1417 net217 net521 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__mux2_1
X_11280_ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__inv_2
XANTENNA__08162__X _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ net225 net1812 net382 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10344__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A2 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ net1710 net222 net526 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1006 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
Xfanout1026 net1030 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
X_10093_ net228 net2262 net388 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07149__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1061 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_184_Left_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ clknet_leaf_60_clk _01375_ net1104 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09153__B _04169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12803_ clknet_leaf_35_clk _00349_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13783_ clknet_leaf_64_clk _01308_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10995_ net907 _05005_ _05015_ net865 vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_54_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12734_ clknet_leaf_39_clk _00280_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__Y _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06675__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12665_ clknet_leaf_58_clk _00211_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10519__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11616_ _05475_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__or2_2
X_12596_ clknet_leaf_96_clk _00142_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11547_ _05404_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__nor2_1
Xhold509 top.DUT.register\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output98_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11478_ _01392_ _05330_ _05305_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13217_ clknet_leaf_41_clk _00763_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10429_ net1933 net237 net512 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07388__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07927__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ clknet_leaf_16_clk _00694_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13079_ clknet_leaf_112_clk _00625_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1209 top.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_183_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08888__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07640_ _02750_ _02752_ _02754_ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__or4_1
XFILLER_0_189_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13492__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07571_ net829 net331 _02669_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__o21a_1
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08104__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09310_ _04339_ _04340_ _04338_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a21o_1
X_06522_ _01630_ _01635_ _01638_ net400 net856 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ _04285_ _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__or2_1
X_06453_ net810 _01535_ net808 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__and3_1
XANTENNA__06666__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09172_ top.pc\[2\] _04209_ _04223_ net873 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a211o_1
X_06384_ top.pad.button_control.r_counter\[14\] top.pad.button_control.r_counter\[13\]
+ top.pad.button_control.r_counter\[12\] top.pad.button_control.r_counter\[11\] vssd1
+ vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__or4_1
XFILLER_0_113_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__C_N top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09604__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08123_ top.DUT.register\[5\]\[16\] net540 _03237_ _03239_ vssd1 vssd1 vccd1 vccd1
+ _03240_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout217_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ top.DUT.register\[8\]\[23\] net556 net544 top.DUT.register\[24\]\[23\] _03170_
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a221o_1
XANTENNA__07091__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07005_ top.DUT.register\[30\]\[19\] net760 net711 top.DUT.register\[25\]\[19\] _02121_
+ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a221o_1
XANTENNA__10164__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07379__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11175__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__A2 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08956_ net1301 net860 net838 _04043_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07907_ top.DUT.register\[4\]\[24\] net551 net657 top.DUT.register\[28\]\[24\] _03023_
+ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ _03955_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout753_A _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ _01878_ _02952_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07769_ top.DUT.register\[11\]\[30\] net702 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ net151 net1830 net372 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06657__A2 _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ _02153_ _04460_ _04463_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a21o_1
XANTENNA__10339__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12450_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[13\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_191_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ top.a1.dataIn\[29\] top.a1.dataIn\[30\] _05231_ vssd1 vssd1 vccd1 vccd1 _05262_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12381_ _06155_ _06156_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__nor2_1
XANTENNA__08803__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _05194_ _05196_ _05198_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10074__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _05131_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07909__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ clknet_leaf_118_clk _00548_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10214_ net154 net2084 net438 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ net865 _05095_ top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__o21a_1
X_10145_ net155 net1864 net442 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_192_Left_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10802__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06593__A1 _01709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07790__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ net160 net1533 net448 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
XANTENNA__12302__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06300__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13835_ clknet_leaf_42_clk _01358_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13766_ clknet_leaf_66_clk _01291_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08508__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ net2000 net151 net484 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XANTENNA__09834__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ clknet_leaf_114_clk _00263_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06648__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ clknet_leaf_61_clk _01230_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__B _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ clknet_leaf_24_clk _00194_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12579_ clknet_leaf_29_clk _00125_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07073__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 top.DUT.register\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold317 top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top.DUT.register\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold339 top.DUT.register\[6\]\[20\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06820__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 _01536_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_2
Xfanout819 _04170_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_2
X_08810_ net398 _03179_ _03180_ net477 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09770__A1 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _04784_ _04789_ _04192_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a21o_1
XANTENNA__07781__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 top.DUT.register\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09074__A _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 top.DUT.register\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net903 top.pc\[19\] net538 _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1028 top.DUT.register\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1039 top.DUT.register\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10668__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ _02523_ _03762_ _03772_ net473 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ net829 _02739_ net468 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09839__B1_N _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_166_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__B _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ top.DUT.register\[19\]\[9\] net673 net641 top.DUT.register\[9\]\[9\] _02670_
+ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_196_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09825__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06505_ _01388_ _01596_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nor2_1
X_07485_ top.DUT.register\[7\]\[7\] net574 net645 top.DUT.register\[10\]\[7\] _02601_
+ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a221o_1
XANTENNA__06639__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ _04261_ _04272_ _04271_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__a21oi_1
X_06436_ top.a1.instruction\[19\] net830 _01552_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__and3b_4
XFILLER_0_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12555__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ net855 _04204_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__and3_2
X_06367_ top.a1.instruction\[13\] top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ _01490_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08106_ top.DUT.register\[6\]\[22\] net577 net684 top.DUT.register\[2\]\[22\] _03222_
+ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a221o_1
XANTENNA__07064__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09086_ _04007_ _04030_ _04072_ _04050_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or4b_1
X_06298_ top.ramload\[24\] net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ _02132_ _03152_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__nor2_1
XANTENNA__06811__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold840 top.DUT.register\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold851 top.DUT.register\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 top.DUT.register\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 top.DUT.register\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 top.DUT.register\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 top.DUT.register\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10622__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net233 net1887 net452 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__mux2_1
XANTENNA__07772__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ net298 net358 _03343_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _05808_ _05809_ _05799_ _05803_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_106_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ net1837 net197 net407 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06878__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _01398_ net127 _05699_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a21o_1
X_13620_ clknet_leaf_92_clk net1158 net996 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
X_10832_ net1945 net208 net493 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11084__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ clknet_leaf_21_clk _01097_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10069__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ net221 net1914 net371 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ clknet_leaf_76_clk _00049_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13482_ clknet_leaf_118_clk _01028_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10694_ net1775 net234 net499 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12433_ clknet_leaf_78_clk top.ru.next_FetchedData\[28\] net1081 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07055__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12364_ net2308 _06143_ _06145_ net814 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _05129_ _05149_ _05161_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12295_ net1206 _06101_ _06103_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08998__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11246_ net872 _05110_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10532__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__B _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ net925 net1364 _01440_ _05088_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a31o_1
X_10128_ net225 net1851 net442 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13084__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10059_ net229 net1575 net448 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XANTENNA__07515__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A3 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06869__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ clknet_leaf_71_clk _01343_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13749_ clknet_leaf_62_clk _01274_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ top.DUT.register\[27\]\[3\] net773 net753 top.DUT.register\[17\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07294__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06221_ _01429_ _01430_ _01434_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[3\] sky130_fd_sc_hd__or3_1
XFILLER_0_170_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10707__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07046__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 top.a1.row1\[2\] vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold114 top.a1.row1\[16\] vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _01164_ vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold136 top.ramaddr\[4\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 top.DUT.register\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _04898_ _04899_ _04897_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o21ai_1
Xhold169 top.DUT.register\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net607 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09743__A1 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _04727_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_4
XANTENNA__10442__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_8
X_09842_ _04836_ _04837_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__and2_1
Xfanout638 _01701_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout649 _01696_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07754__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ top.a1.dataIn\[10\] _04766_ _04769_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_
+ sky130_fd_sc_hd__a211o_1
X_06985_ top.DUT.register\[1\]\[20\] net781 net711 top.DUT.register\[25\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout284_A _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _03106_ _03802_ _02153_ _03103_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_198_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10949__Y _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08655_ _02517_ _03748_ _03756_ net467 _03754_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout451_A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ top.DUT.register\[11\]\[11\] net700 net644 top.DUT.register\[10\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
X_08586_ _02824_ _03690_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__or2_1
XANTENNA__11066__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07537_ top.DUT.register\[20\]\[13\] net560 net667 top.DUT.register\[31\]\[13\] _02653_
+ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a221o_1
XANTENNA__07809__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07987__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07285__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _02578_ _02580_ _02582_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__or4_1
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09207_ top.pc\[5\] _01808_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06419_ top.a1.instruction\[17\] top.a1.instruction\[18\] net830 vssd1 vssd1 vccd1
+ vccd1 _01536_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10617__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ _01735_ _01744_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__nor2_1
XANTENNA__08234__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ net913 _01595_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor2_2
XFILLER_0_121_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09069_ _03574_ _03618_ _04121_ _03598_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ net82 net880 net848 net1256 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a22o_1
XANTENNA__07993__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _05915_ _05921_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 top.DUT.register\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 top.DUT.register\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold692 top.DUT.register\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ top.a1.dataInTemp\[9\] net798 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__or2_1
XANTENNA__10352__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_102_clk _00528_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09442__A _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _05790_ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09161__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11864_ _05707_ net128 vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ clknet_leaf_55_clk _01144_ net1097 vssd1 vssd1 vccd1 vccd1 top.ramload\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_45_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10815_ net146 net1844 net413 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ _01397_ net129 _05625_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ clknet_leaf_38_clk _01080_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10746_ net157 net1819 net414 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XANTENNA__07276__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08473__B2 _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ clknet_leaf_56_clk _01011_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10527__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10677_ net168 net1556 net421 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12416_ clknet_leaf_54_clk top.ru.next_FetchedData\[11\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07028__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ clknet_leaf_99_clk _00942_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09973__A1 _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ top.pad.button_control.r_counter\[0\] net1250 _06134_ vssd1 vssd1 vccd1 vccd1
+ _01354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12278_ net1182 _06091_ net1117 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09725__A1 top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ net871 _05015_ _05029_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__and3_1
XANTENNA__10262__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06770_ top.DUT.register\[9\]\[29\] net715 net754 top.DUT.register\[18\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08667__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__A _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__Y _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _03523_ _02837_ _02587_ _02468_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _03411_ _03483_ net314 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ top.DUT.register\[15\]\[7\] net806 net803 top.DUT.register\[31\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XANTENNA__07267__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08255__X _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07600__A _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07253_ net286 _02368_ _02369_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10437__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06204_ top.a1.halfData\[1\] top.a1.halfData\[2\] top.a1.halfData\[3\] vssd1 vssd1
+ vccd1 vccd1 _01424_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07019__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ top.DUT.register\[30\]\[11\] net761 _02287_ _02300_ vssd1 vssd1 vccd1 vccd1
+ _02301_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09413__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09527__A _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _05114_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _04998_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10172__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_8
Xfanout435 _04980_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
Xfanout446 _04967_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _03781_ net454 net533 _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__o211a_2
Xfanout457 _04736_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
Xfanout468 _02618_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_4
Xfanout479 _05263_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10900__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ net237 top.DUT.register\[1\]\[7\] net392 vssd1 vssd1 vccd1 vccd1 _00129_
+ sky130_fd_sc_hd__mux2_1
X_06968_ top.DUT.register\[29\]\[21\] net785 net720 top.DUT.register\[26\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a22o_1
XANTENNA__06886__A _01993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _03107_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__or2_1
X_09687_ _04697_ _04700_ _04704_ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__or4_1
XFILLER_0_179_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ top.DUT.register\[6\]\[24\] net599 net773 top.DUT.register\[27\]\[24\] _02015_
+ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _03717_ _02641_ _02638_ _02244_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net301 _03472_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10600_ net214 net2130 net422 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ top.a1.dataIn\[14\] _05386_ _05401_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06466__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ net223 net2112 net426 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10347__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ clknet_leaf_10_clk _00796_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10462_ net237 net2171 net508 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12201_ _06053_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__and2_1
XANTENNA__11481__A1_N top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ clknet_leaf_120_clk _00727_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10393_ net2021 net252 net515 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12132_ _05953_ _05986_ _05990_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12063_ _05919_ _05920_ _05923_ _05892_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a22o_2
XANTENNA__09156__B _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net864 _05029_ _05030_ net869 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1
+ _05031_ sky130_fd_sc_hd__a32o_1
Xfanout980 net982 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10810__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08487__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ clknet_leaf_46_clk _00511_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11916_ _05743_ _05761_ _05774_ _05775_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07404__B _01733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08694__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ clknet_leaf_14_clk _00442_ net981 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11847_ _05693_ _05690_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11778_ _05604_ _05632_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13517_ clknet_leaf_113_clk _01063_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06457__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10729_ net226 net2236 net414 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10257__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload12 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinvlp_4
X_13448_ clknet_leaf_31_clk _00994_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload23 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__bufinv_16
Xclkload45 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload56 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_16
X_13379_ clknet_leaf_34_clk _00925_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload67 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinv_2
Xclkload78 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_4
XANTENNA__07957__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload89 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__inv_8
XFILLER_0_140_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08251__A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_11__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _02003_ _03053_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__or2_1
XFILLER_0_208_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07871_ top.DUT.register\[28\]\[27\] net655 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_79_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08382__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ _04633_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ _01934_ _01936_ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__or3_1
XANTENNA__10720__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _04569_ _04570_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06753_ top.DUT.register\[7\]\[28\] net708 net755 top.DUT.register\[18\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09472_ _04504_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07488__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06684_ _01738_ net285 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ net281 _03533_ _03531_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06696__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_A _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08354_ _02552_ _03442_ _02558_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a21o_1
XANTENNA__08437__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07305_ top.DUT.register\[21\]\[1\] net611 net591 top.DUT.register\[20\]\[1\] _02421_
+ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10167__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload6 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_8
X_08285_ _03397_ _03399_ net287 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_2
XFILLER_0_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout414_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ top.DUT.register\[6\]\[8\] net598 net594 top.DUT.register\[8\]\[8\] _02352_
+ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a221o_1
XANTENNA__07660__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07167_ net348 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__inv_2
X_07098_ top.DUT.register\[8\]\[15\] net594 net772 top.DUT.register\[27\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout783_A _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout221 _04781_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 _04772_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 _04742_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_208_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 net256 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_2
Xfanout265 _04750_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_2
Xfanout276 _01858_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
X_09808_ _04410_ net362 _04806_ _04769_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a211o_1
XANTENNA__10630__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
X_09739_ _03465_ net456 net536 _04749_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__o211a_4
XFILLER_0_202_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08125__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12750_ clknet_leaf_95_clk _00296_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07479__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11701_ _05558_ _05561_ _05556_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12681_ clknet_leaf_26_clk _00227_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08428__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11632_ _05424_ _05460_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_194_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08428__B2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10077__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ _05417_ _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ clknet_leaf_103_clk _00848_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10514_ net158 net2033 net379 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__mux2_1
X_11494_ _05325_ _05326_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13233_ clknet_leaf_9_clk _00779_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net1516 net172 net510 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
XANTENNA__10805__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07403__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13164_ clknet_leaf_3_clk _00710_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10376_ net1665 net179 net431 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
X_12115_ _05953_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13095_ clknet_leaf_49_clk _00641_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12046_ _05884_ _05895_ _05904_ _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__a22o_1
XANTENNA__12839__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08116__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12421__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ clknet_leaf_104_clk _00494_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09864__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12879_ clknet_leaf_21_clk _00425_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08070_ top.DUT.register\[21\]\[17\] net569 net565 top.DUT.register\[23\]\[17\] _03186_
+ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a221o_1
Xclkload101 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__07642__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ top.DUT.register\[27\]\[18\] net770 _02137_ vssd1 vssd1 vccd1 vccd1 _02138_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06850__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10715__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06401__A_N top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__A1 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ net461 _04045_ _04058_ net465 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__o22a_1
XFILLER_0_87_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07923_ top.DUT.register\[6\]\[25\] net579 net686 top.DUT.register\[2\]\[25\] _03039_
+ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a221o_1
Xhold18 top.ramstore\[0\] vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 top.a1.data\[1\] vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10450__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ top.DUT.register\[7\]\[26\] net574 net645 top.DUT.register\[10\]\[26\] _02970_
+ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__a221o_1
X_06805_ top.DUT.register\[28\]\[31\] net740 net594 top.DUT.register\[8\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07785_ _01920_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__or2_1
XFILLER_0_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08107__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ net137 _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_203_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06736_ _01843_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_203_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08658__B2 _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06669__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ top.pc\[20\] _04477_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__or2_1
X_06667_ top.DUT.register\[1\]\[1\] net705 _01783_ vssd1 vssd1 vccd1 vccd1 _01784_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout629_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08406_ _02560_ _03489_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__and2b_1
XANTENNA__07331__Y _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09386_ net854 _01803_ net619 _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__o22a_4
XANTENNA__07881__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06598_ top.a1.instruction\[24\] top.a1.instruction\[25\] top.a1.instruction\[26\]
+ top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08337_ _01775_ _03449_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nor2_1
XANTENNA__09083__A1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07094__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ net1340 _01511_ net838 _03383_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a22o_1
XANTENNA__07633__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06841__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ top.DUT.register\[4\]\[9\] net582 net757 top.DUT.register\[3\]\[9\] _02335_
+ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a221o_1
XANTENNA__10625__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ net297 net339 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Right_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10230_ net230 net2062 net384 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ net1455 net226 net525 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1019 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_2
Xfanout1027 net1030 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
Xfanout1038 net1050 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
X_10092_ net232 net1916 net388 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_2
XFILLER_0_199_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10360__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09434__B _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13851_ clknet_leaf_60_clk _01374_ net1104 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12802_ clknet_leaf_12_clk _00348_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13782_ clknet_leaf_65_clk _01307_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10994_ top.a1.dataInTemp\[0\] _05009_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ clknet_leaf_120_clk _00279_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12664_ clknet_leaf_37_clk _00210_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07872__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11615_ _05443_ net207 _05447_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10883__X _05001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ clknet_leaf_109_clk _00141_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _05388_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06832__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10535__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _01392_ _05330_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ clknet_leaf_13_clk _00762_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ net1669 net246 net511 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13147_ clknet_leaf_5_clk _00693_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10359_ net1538 net254 net433 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ clknet_leaf_102_clk _00624_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _05888_ _05889_ _05858_ _05864_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10270__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire332_A _02687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06899__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07570_ _02671_ _02673_ _02677_ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__nor4_2
XTAP_TAPCELL_ROW_66_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07432__X _02549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ _01637_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09240_ _04286_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
X_06452_ net810 _01527_ net808 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ net916 net910 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nand2_2
X_06383_ net1977 _01500_ top.ru.next_read_i vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__o21a_1
XANTENNA__13674__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07076__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ top.DUT.register\[22\]\[16\] net552 net655 top.DUT.register\[28\]\[16\] _03238_
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07615__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ top.DUT.register\[2\]\[23\] net683 net655 top.DUT.register\[28\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a22o_1
XANTENNA__10445__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ top.DUT.register\[27\]\[19\] net770 net766 top.DUT.register\[11\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1021_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ net904 top.pc\[29\] net538 _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ top.DUT.register\[30\]\[24\] net697 net673 top.DUT.register\[19\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_1
XANTENNA__10180__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ net461 _03960_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07000__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__C top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _01878_ _02952_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A1 top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07768_ top.DUT.register\[4\]\[30\] net551 net629 top.DUT.register\[29\]\[30\] _02884_
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _04519_ _04520_ _04521_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o21ai_2
X_06719_ top.DUT.register\[10\]\[3\] net646 net625 top.DUT.register\[16\]\[3\] _01835_
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07699_ top.DUT.register\[22\]\[12\] net552 net635 top.DUT.register\[25\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ _04472_ _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07854__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ net841 _01750_ net619 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11400_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__inv_2
XANTENNA__07067__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ net1789 _06153_ net815 vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07606__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ top.a1.row2\[27\] _05134_ _05140_ top.a1.row1\[59\] _05142_ vssd1 vssd1 vccd1
+ vccd1 _05199_ sky130_fd_sc_hd__a221o_1
XANTENNA__06814__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11262_ top.lcd.nextState\[1\] _01382_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13001_ clknet_leaf_26_clk _00547_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10213_ net158 net2234 net440 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
X_11193_ net1688 _05099_ _05096_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
XANTENNA__08031__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10144_ net159 net1667 net443 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10090__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ net162 net1813 net449 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ clknet_leaf_42_clk _01357_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13765_ clknet_leaf_66_clk _01290_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ net1392 net154 net481 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XANTENNA__08098__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08508__B _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12716_ clknet_leaf_3_clk _00262_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_13696_ clknet_leaf_61_clk _01229_ net1110 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07845__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ clknet_leaf_49_clk _00193_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12578_ clknet_leaf_10_clk _00124_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06805__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10265__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11529_ _05363_ _05364_ _05346_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 top.DUT.register\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 top.DUT.register\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 top.DUT.register\[31\]\[0\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_185_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08022__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout809 _01517_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09770__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1007 top.DUT.register\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07146__Y _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ net461 _03823_ _03837_ net466 _03835_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1018 top.DUT.register\[17\]\[17\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 top.DUT.register\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ net271 _03595_ _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07622_ _02729_ _02738_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nor2_4
XFILLER_0_177_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_200_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07553_ top.DUT.register\[30\]\[9\] net697 net645 top.DUT.register\[10\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06504_ net914 _01491_ _01484_ top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01621_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_196_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07297__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ top.DUT.register\[30\]\[7\] net697 net629 top.DUT.register\[29\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_200_Right_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _02489_ _02529_ _04260_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a21o_1
X_06435_ top.a1.instruction\[15\] top.a1.instruction\[16\] _01528_ vssd1 vssd1 vccd1
+ vccd1 _01552_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1069_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ _04169_ _04201_ _04205_ _04078_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__o221a_1
X_06366_ net912 top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08105_ top.DUT.register\[18\]\[22\] net660 net656 top.DUT.register\[28\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a22o_1
XANTENNA__10175__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ _03637_ _03664_ _04136_ _04137_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_15_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06297_ net1241 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[23\] sky130_fd_sc_hd__and2_1
XFILLER_0_114_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08036_ _02132_ _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold830 top.DUT.register\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 top.DUT.register\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold852 top.DUT.register\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout696_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 top.DUT.register\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A1 _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 top.DUT.register\[10\]\[13\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10903__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 top.DUT.register\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 top.DUT.register\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07221__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net238 net1983 net452 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout863_A _05053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net306 _03705_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08869_ _02982_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10900_ net1502 net201 net406 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11880_ _01398_ _05699_ net127 vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nand3_1
XFILLER_0_168_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ top.DUT.register\[27\]\[13\] net212 net493 vssd1 vssd1 vccd1 vccd1 _00967_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13550_ clknet_leaf_97_clk _01096_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07288__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ net223 net2268 net370 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07827__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12501_ clknet_leaf_88_clk _00048_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13481_ clknet_leaf_26_clk _01027_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09029__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ net1347 net236 net499 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ clknet_leaf_78_clk top.ru.next_FetchedData\[27\] net1081 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[27\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_33_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ top.pad.button_control.r_counter\[7\] _06143_ vssd1 vssd1 vccd1 vccd1 _06145_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10085__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08063__B _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11314_ net900 _05148_ _05143_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_200_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09727__X _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07460__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12294_ net1206 _06101_ net1118 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11245_ net1856 net403 _04682_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08004__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07212__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ net64 net884 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__and2_1
XANTENNA__13693__Q top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ net231 net1638 net444 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_42_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ net234 net1598 net448 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06738__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13817_ clknet_leaf_72_clk _01342_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07279__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13748_ clknet_leaf_67_clk _01273_ vssd1 vssd1 vccd1 vccd1 top.lcd.lcd_rs sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07818__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_88_clk _01220_ net1018 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06220_ top.a1.hexop\[2\] top.a1.hexop\[1\] top.a1.hexop\[3\] top.a1.hexop\[4\] vssd1
+ vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08254__A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 top.a1.row1\[123\] vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 top.DUT.register\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold137 net85 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 top.ramstore\[31\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__C1 _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold159 top.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ top.pc\[25\] _04576_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nor2_1
XANTENNA__10723__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ _04824_ _04825_ _04826_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__o21a_1
Xfanout617 _04727_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09743__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout628 net630 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06557__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 _01699_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_8
X_09772_ net818 _04322_ net816 top.pc\[10\] vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__a2bb2o_1
X_06984_ top.DUT.register\[2\]\[20\] net775 _02100_ vssd1 vssd1 vccd1 vccd1 _02101_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08723_ net1331 net859 net837 _03821_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_198_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ _02720_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ top.DUT.register\[3\]\[11\] net692 net549 top.DUT.register\[4\]\[11\] _02721_
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a221o_1
X_08585_ _03640_ _03689_ _02741_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ top.DUT.register\[6\]\[13\] net576 net679 top.DUT.register\[26\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
XANTENNA__07809__A2 _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ top.DUT.register\[8\]\[6\] net558 net637 top.DUT.register\[25\]\[6\] _02583_
+ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a221o_1
XANTENNA__08482__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09206_ _04254_ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06418_ top.a1.instruction\[15\] top.a1.instruction\[16\] net830 vssd1 vssd1 vccd1
+ vccd1 _01535_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07690__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ net312 _02201_ net271 _02371_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__o221a_1
XANTENNA__08164__A _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09137_ top.a1.instruction\[11\] _04181_ _04182_ _04189_ vssd1 vssd1 vccd1 vccd1
+ _04190_ sky130_fd_sc_hd__and4_2
X_06349_ _01332_ _01333_ _01468_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__and3b_1
XFILLER_0_20_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _03355_ _03403_ _03439_ net277 vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout980_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06796__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ top.DUT.register\[23\]\[19\] net565 net631 top.DUT.register\[27\]\[19\] _03135_
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a221o_1
XANTENNA__10633__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold660 top.DUT.register\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 top.DUT.register\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net1181 _05042_ net480 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
Xhold682 top.DUT.register\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 top.DUT.register\[28\]\[22\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06548__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_101_clk _00527_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11932_ _05764_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09442__B _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__A1 _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ _05717_ _05722_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06720__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11057__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ clknet_leaf_53_clk _01143_ net1075 vssd1 vssd1 vccd1 vccd1 top.ramload\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10814_ net147 net2127 net410 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11794_ _01397_ _05625_ net129 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ clknet_leaf_120_clk _01079_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ net159 net1809 net415 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XANTENNA__09670__A1 _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10808__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13464_ clknet_leaf_33_clk _01010_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10676_ net170 top.DUT.register\[22\]\[23\] net418 vssd1 vssd1 vccd1 vccd1 _00817_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12308__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12415_ clknet_leaf_55_clk top.ru.next_FetchedData\[10\] net1097 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12446__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ clknet_leaf_111_clk _00941_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12346_ top.pad.button_control.r_counter\[0\] net1250 net815 vssd1 vssd1 vccd1 vccd1
+ _06134_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06787__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12277_ _06091_ _06092_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10543__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ net908 net909 _05095_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ net923 net1281 net875 _05079_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09352__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11048__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ net342 net334 net321 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux2_1
XANTENNA__06992__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07321_ _02431_ _02433_ _02435_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__or4_4
XFILLER_0_46_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07252_ net291 _02286_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07672__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06203_ top.a1.halfData\[3\] _01422_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__nand2_1
XANTENNA__11122__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ top.DUT.register\[6\]\[11\] net597 net708 top.DUT.register\[7\]\[11\] _02299_
+ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a221o_1
XANTENNA__09413__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07424__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06778__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10453__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09527__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _05114_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06232__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 net417 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_6
Xfanout425 _04992_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_8
Xfanout436 _04980_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_6
XFILLER_0_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _04821_ _04819_ _04818_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__or3b_1
Xfanout447 _04967_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
Xfanout458 net460 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 net471 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
X_06967_ top.DUT.register\[6\]\[21\] net597 net761 top.DUT.register\[30\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a22o_1
X_09755_ _03581_ net456 net535 _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout561_A _01673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__B _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _03777_ _03804_ _03205_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09686_ _04699_ _04703_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ top.DUT.register\[16\]\[24\] net724 net762 top.DUT.register\[30\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ net1326 net858 net836 _03739_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1091_X net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ net271 _03470_ _03478_ net274 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ _02629_ _02631_ _02633_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08499_ net277 _03310_ _03341_ net270 vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__a22o_1
XANTENNA__10628__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10530_ net228 net2039 net428 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07663__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10461_ net247 net2176 net508 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12200_ _06052_ _06054_ _06049_ _06050_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07415__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ clknet_leaf_18_clk _00726_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10392_ net2010 net253 net515 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__mux2_1
XANTENNA__06769__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ _05975_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nor2_1
XANTENNA__10363__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12062_ _05867_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__nand2_1
Xhold490 top.DUT.register\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ top.a1.dataInTemp\[4\] net798 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or2_1
XANTENNA__07194__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net978 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_2
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06941__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12964_ clknet_leaf_29_clk _00510_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1190 top.DUT.register\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ _05774_ _05775_ _05743_ _05761_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_142_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_32_clk _00441_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12227__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11846_ _05703_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _05605_ _05634_ _05635_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__nand4_1
XANTENNA__10538__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13516_ clknet_leaf_115_clk _01062_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10728_ net231 net2032 net416 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13447_ clknet_leaf_56_clk _00993_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10659_ net245 net1557 net420 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__mux2_1
Xclkload13 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_51_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload24 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload35 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_12
XFILLER_0_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload46 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_58_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09946__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_11_clk _00924_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload57 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_12
Xclkload68 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_8
Xclkload79 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_16
X_12329_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__inv_2
XANTENNA__10273__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ top.DUT.register\[3\]\[27\] net691 net651 top.DUT.register\[17\]\[27\] _02986_
+ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a221o_1
XANTENNA__07185__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ top.DUT.register\[24\]\[31\] net587 net713 top.DUT.register\[25\]\[31\] _01937_
+ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a221o_1
XANTENNA__08382__B2 _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09540_ top.pc\[25\] _04557_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__and2_1
X_06752_ top.DUT.register\[25\]\[28\] net713 net759 top.DUT.register\[2\]\[28\] _01868_
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ top.pc\[21\] _04494_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06683_ net313 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08422_ _03352_ _03402_ _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__and3b_1
XANTENNA__12218__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__B _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__X _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08353_ net1462 net861 net838 _03466_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10448__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout142_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ top.DUT.register\[3\]\[1\] net783 net733 top.DUT.register\[23\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08284_ net319 _01942_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__nand2_1
XANTENNA__07645__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload7 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06999__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07235_ top.DUT.register\[1\]\[8\] net780 net772 top.DUT.register\[27\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1051_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ _02267_ _02277_ _02280_ _02282_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__nor4_2
XANTENNA__09538__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08070__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ top.DUT.register\[17\]\[15\] net776 _02213_ vssd1 vssd1 vccd1 vccd1 _02214_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06233__Y _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09825__X _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__A _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 _04823_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 _04805_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout776_A _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 _04781_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_1
Xfanout233 _04772_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10911__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout244 net247 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_208_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07176__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _04750_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_1
XANTENNA__08606__A1_N net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__B2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_2
X_09807_ net818 _04417_ _04766_ top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _04806_
+ sky130_fd_sc_hd__a2bb2o_1
Xfanout288 _01775_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ _03109_ _03111_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__or3_1
XFILLER_0_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06923__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09738_ top.a1.dataIn\[3\] _01499_ _04736_ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_2_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net909 _04687_ _04690_ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__o21a_1
XFILLER_0_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ _05524_ _05559_ _05523_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__nor3b_1
XANTENNA__06687__A1 top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ clknet_leaf_26_clk _00226_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06687__B2 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11631_ _05462_ _05490_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12720__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11043__A _01400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07636__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ _05395_ _05396_ net248 _05397_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07100__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ net162 net1377 net381 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13301_ clknet_leaf_82_clk _00847_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11493_ _05334_ _05337_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__nor3_1
X_13232_ clknet_leaf_116_clk _00778_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10444_ net1676 net177 net510 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08061__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ clknet_leaf_4_clk _00709_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10093__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10375_ net1610 net183 net431 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _05945_ _05955_ _05946_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__a21o_1
XANTENNA__09735__X _04747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13094_ clknet_leaf_47_clk _00640_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ _05888_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_53_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12321__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12947_ clknet_leaf_108_clk _00493_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__Y _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12878_ clknet_leaf_95_clk _00424_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ _05653_ _05688_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__xor2_2
XANTENNA__10268__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload102 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_8
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07020_ top.DUT.register\[6\]\[18\] net596 net715 top.DUT.register\[9\]\[18\] _02136_
+ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_188_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08052__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08971_ _02905_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__xnor2_1
X_07922_ top.DUT.register\[30\]\[25\] net698 net571 top.DUT.register\[21\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a22o_1
XANTENNA__10731__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 _01161_ vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ top.DUT.register\[20\]\[26\] net562 net649 top.DUT.register\[12\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a22o_1
X_06804_ net324 _01919_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__nand2_1
X_07784_ net828 _02900_ _02618_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13879__1139 vssd1 vssd1 vccd1 vccd1 _13879__1139/HI net1139 sky130_fd_sc_hd__conb_1
X_06735_ _01845_ _01847_ _01849_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__or4_1
XANTENNA__09821__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12549__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09523_ _04550_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_203_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09855__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1099_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ top.pc\[20\] _04477_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06666_ top.DUT.register\[14\]\[1\] net665 net638 top.DUT.register\[25\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09540__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08405_ net469 _03505_ _03516_ _02522_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10178__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _01595_ _01805_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06597_ top.a1.instruction\[28\] top.a1.instruction\[29\] top.a1.instruction\[30\]
+ top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout524_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09967__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08336_ _03449_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07618__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08267_ net905 top.pc\[1\] net539 _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10906__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07218_ top.DUT.register\[8\]\[9\] net594 net762 top.DUT.register\[30\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a22o_1
XANTENNA__09268__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08198_ net321 _02428_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08043__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ top.DUT.register\[16\]\[12\] net725 net711 top.DUT.register\[25\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09791__B1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net1507 net228 net526 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1021 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10641__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
X_10091_ net236 net1732 net388 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
Xfanout1028 net1030 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07149__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1039 net1041 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13850_ clknet_leaf_59_clk _01373_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12801_ clknet_leaf_43_clk _00347_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10993_ net907 _05008_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__or2_1
X_13781_ clknet_leaf_65_clk _01306_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ clknet_leaf_17_clk _00278_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07857__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09116__C_N _04168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__Y _05053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10088__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ clknet_leaf_107_clk _00209_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08066__B _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07609__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ _05443_ _05447_ net207 vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__and3_1
X_12594_ clknet_leaf_106_clk _00140_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11545_ _05387_ net248 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__nand2_1
XANTENNA__10816__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ _05314_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__xor2_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10427_ net1463 net249 net511 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
X_13215_ clknet_leaf_22_clk _00761_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07388__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10358_ net2284 net268 net432 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ clknet_leaf_15_clk _00692_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10551__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ clknet_leaf_100_clk _00623_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10289_ net2181 net263 net524 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__mux2_1
XANTENNA__06601__Y _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _05804_ _05854_ _05839_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_183_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08888__A2 _03977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_clk_X clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06520_ top.a1.instruction\[21\] _01634_ _01636_ vssd1 vssd1 vccd1 vccd1 _01637_
+ sky130_fd_sc_hd__a21oi_2
XANTENNA__07848__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06451_ top.a1.instruction\[15\] top.a1.instruction\[16\] net810 _01520_ vssd1 vssd1
+ vccd1 vccd1 _01568_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09787__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ _04091_ net138 _04218_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06382_ _01501_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ top.DUT.register\[15\]\[16\] net687 net631 top.DUT.register\[27\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10726__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08052_ top.DUT.register\[15\]\[23\] net687 net643 top.DUT.register\[10\]\[23\] _03168_
+ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07003_ top.DUT.register\[14\]\[19\] net792 net604 top.DUT.register\[22\]\[19\] _02119_
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08025__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07379__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09773__B1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10461__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _04040_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ top.DUT.register\[7\]\[24\] net575 net682 top.DUT.register\[26\]\[24\] _03021_
+ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_90_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08885_ net465 _03965_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11883__A1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07767_ top.DUT.register\[31\]\[30\] net669 net666 top.DUT.register\[14\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a22o_1
XANTENNA__09289__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout739_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09506_ _04536_ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nand2b_1
X_06718_ top.DUT.register\[2\]\[3\] net685 net638 top.DUT.register\[25\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07698_ top.DUT.register\[6\]\[12\] net576 net663 top.DUT.register\[14\]\[12\] _02814_
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07303__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09437_ _04454_ _04455_ _04456_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o21ai_1
X_06649_ top.DUT.register\[26\]\[2\] net680 net672 top.DUT.register\[19\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _04394_ _04396_ _04392_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08319_ _02203_ _03429_ _03432_ net274 vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10636__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09299_ top.a1.instruction\[31\] _01640_ net857 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_4_13__f_clk_X clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ top.a1.row1\[107\] _05149_ _05155_ top.a1.row1\[19\] _05197_ vssd1 vssd1
+ vccd1 vccd1 _05198_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _05127_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__nor2_1
XANTENNA__08016__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10212_ net162 net2055 net441 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13000_ clknet_leaf_26_clk _00546_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09764__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _01421_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nor2_1
X_10143_ net164 net1503 net445 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XANTENNA__10371__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09516__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net166 net1807 net449 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
XANTENNA__09461__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ clknet_leaf_42_clk _01356_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06750__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09180__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ clknet_leaf_65_clk _01289_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10976_ net1586 net160 net483 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12715_ clknet_leaf_6_clk _00261_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13695_ clknet_leaf_61_clk _01228_ net1110 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ clknet_leaf_21_clk _00192_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06541__A_N top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10546__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_104_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12577_ clknet_leaf_44_clk _00123_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _05387_ _05388_ _05383_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold308 top.DUT.register\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08007__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 top.DUT.register\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
X_13878__1138 vssd1 vssd1 vccd1 vccd1 _13878__1138/HI net1138 sky130_fd_sc_hd__conb_1
X_11459_ _05289_ _05319_ _05293_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_185_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09755__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ clknet_leaf_27_clk _00675_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10281__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07781__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 top.DUT.register\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 top.DUT.register\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _01802_ _03570_ _03770_ net272 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__o22a_1
XANTENNA__08539__X _03646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07533__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07621_ _02731_ _02733_ _02735_ _02737_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__or4_2
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ net825 _02668_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__or2_1
XANTENNA__13641__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06503_ _01619_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_196_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08494__B1 _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07483_ _02593_ _02595_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ _02468_ _02566_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06434_ net811 _01550_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__nor2_4
XANTENNA__13682__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09153_ _04200_ _04169_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06365_ net912 top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__nor2_1
XANTENNA__10456__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout222_A _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ top.DUT.register\[11\]\[22\] net700 net549 top.DUT.register\[4\]\[22\] _03220_
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _03684_ _03706_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06235__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06296_ net1192 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[22\] sky130_fd_sc_hd__and2_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ net825 _03151_ _02617_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold820 top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08721__Y _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 top.DUT.register\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold842 top.DUT.register\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 top.DUT.register\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold864 top.DUT.register\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 top.DUT.register\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09210__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 top.DUT.register\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 top.DUT.register\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ net244 net1657 net452 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__mux2_1
XANTENNA__07772__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _02932_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__xor2_1
XANTENNA__06980__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__C top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _03056_ _03939_ _03057_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__a21boi_1
XANTENNA__08721__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ top.DUT.register\[30\]\[28\] net697 net570 top.DUT.register\[21\]\[28\] _02935_
+ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06732__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _03858_ _03893_ _03128_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ net1571 net216 net493 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12889__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10761_ net228 net1890 net372 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ clknet_leaf_89_clk _00047_ net1015 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10692_ net2197 net244 net499 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
X_13480_ clknet_leaf_26_clk _01026_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ clknet_leaf_78_clk top.ru.next_FetchedData\[26\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[26\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10366__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12147__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _06143_ _06144_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06799__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11313_ net1213 net843 _05181_ net1115 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ _06101_ _06102_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11244_ _05122_ net1240 net402 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__mux2_1
XANTENNA__09737__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net925 net1996 net877 _05087_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a31o_1
X_10126_ net232 net1787 net444 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XANTENNA__09743__X _04753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_180_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10057_ net239 net2288 net449 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07515__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07704__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06723__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload0_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ clknet_leaf_72_clk _01341_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13747_ clknet_leaf_67_clk _01272_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfxtp_1
X_10959_ net1401 net230 net483 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13678_ clknet_leaf_88_clk _01219_ net1018 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ clknet_leaf_101_clk _00175_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08779__B2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 net116 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _01181_ vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 top.ramstore\[1\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ top.pc\[18\] _04460_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__xnor2_1
Xfanout607 _01533_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_4
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07754__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ net228 net1581 net392 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
X_06983_ top.DUT.register\[15\]\[20\] net805 net801 top.DUT.register\[31\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08722_ net903 top.pc\[18\] net538 _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_198_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _02640_ _03734_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout172_A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07604_ top.DUT.register\[18\]\[11\] net660 net648 top.DUT.register\[12\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a22o_1
X_08584_ _02742_ _02798_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07535_ top.DUT.register\[3\]\[13\] net691 net671 top.DUT.register\[19\]\[13\] _02651_
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1081_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout437_A _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07466_ top.DUT.register\[29\]\[6\] net629 net625 top.DUT.register\[16\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ top.pc\[5\] _04239_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06417_ net811 _01518_ _01528_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__and3_4
XFILLER_0_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _02511_ _02513_ net272 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09975__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06348_ _01334_ _01477_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__and2_1
X_09136_ _01662_ _04184_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and3_1
X_09067_ _03629_ _03666_ _03687_ _03708_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or4bb_1
XANTENNA__10914__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06279_ net1848 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[5\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_116_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ top.DUT.register\[5\]\[19\] net540 net647 top.DUT.register\[12\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a22o_1
XANTENNA__07993__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 top.pad.button_control.r_counter\[13\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 top.DUT.register\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 top.DUT.register\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 top.ramstore\[22\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 top.DUT.register\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _01417_ _04669_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ clknet_leaf_96_clk _00526_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11931_ _05753_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06705__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11862_ _05680_ _05719_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877__1137 vssd1 vssd1 vccd1 vccd1 _13877__1137/HI net1137 sky130_fd_sc_hd__conb_1
XFILLER_0_196_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13601_ clknet_leaf_56_clk _01142_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramload\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ net151 net2104 net412 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__mux2_1
X_11793_ top.a1.dataIn\[8\] net129 vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_45_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ clknet_leaf_51_clk _01078_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ net164 net2290 net416 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07130__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13463_ clknet_leaf_112_clk _01009_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10096__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ net174 net1826 net419 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12414_ clknet_leaf_54_clk top.ru.next_FetchedData\[9\] net1099 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13394_ clknet_leaf_106_clk _00940_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12345_ top.pad.button_control.r_counter\[0\] net815 vssd1 vssd1 vccd1 vccd1 _01353_
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_189_Left_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10824__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12276_ net1715 _06090_ net1117 vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08090__A _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09186__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ net1334 net405 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07197__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ net54 net882 vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06944__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ net164 net2298 net388 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
X_11089_ net102 net885 net849 net1227 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__a22o_1
XANTENNA__07434__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_198_Left_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06992__B _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07320_ top.DUT.register\[3\]\[7\] net783 net586 top.DUT.register\[24\]\[7\] _02436_
+ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07121__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07251_ _02327_ _02367_ net313 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06202_ top.a1.halfData\[2\] top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 _01422_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__09795__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07182_ top.DUT.register\[18\]\[11\] net755 net748 top.DUT.register\[1\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10734__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07975__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__A1_N net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout404 _05107_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
XANTENNA__06232__B net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 net417 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_4
Xfanout426 net429 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
Xfanout437 _04980_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09824__A _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _04425_ net362 net329 top.a1.dataIn\[16\] net364 vssd1 vssd1 vccd1 vccd1
+ _04821_ sky130_fd_sc_hd__a221o_1
Xfanout448 _04967_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_6
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06935__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ top.pc\[7\] net817 net457 _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a211o_1
X_06966_ top.DUT.register\[25\]\[21\] net712 _02080_ _02082_ vssd1 vssd1 vccd1 vccd1
+ _02083_ sky130_fd_sc_hd__a211o_1
X_08705_ _03204_ _03253_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09685_ _04691_ _04701_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
X_06897_ top.DUT.register\[15\]\[24\] net806 net802 top.DUT.register\[31\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net902 top.pc\[14\] net537 _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__a22o_1
XANTENNA__07360__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10909__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _02824_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09637__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_202_Left_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout819_A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ top.DUT.register\[21\]\[14\] net568 net564 top.DUT.register\[23\]\[14\] _02634_
+ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07112__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ _02695_ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06466__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ top.a1.instruction\[27\] net857 _01615_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__A_N _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ net249 net1658 net508 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ _01514_ _01604_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nor2_1
XANTENNA__10644__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ net1490 net268 net516 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08612__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12130_ _05972_ _05985_ _05953_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06423__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Left_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _05885_ _05887_ _05891_ _05894_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a31o_1
Xhold480 top.DUT.register\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 top.ramstore\[25\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ top.a1.data\[0\] net797 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__or2_1
XANTENNA__06926__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net1021 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
Xfanout971 net978 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
Xfanout982 net994 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13714__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ clknet_leaf_34_clk _00509_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_84_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1180 top.DUT.register\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 top.DUT.register\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11914_ top.a1.dataIn\[5\] _05699_ _05740_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__or3_1
X_12894_ clknet_leaf_37_clk _00440_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11845_ _05704_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__and2_1
XFILLER_0_185_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10819__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11776_ _05596_ _05636_ _05632_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07103__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ clknet_leaf_12_clk _01061_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06457__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10727_ net232 net1648 net416 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13446_ clknet_leaf_45_clk _00992_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10658_ net252 net1794 net420 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08372__X _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload14 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_8
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload25 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__bufinv_16
Xclkload36 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10554__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ clknet_leaf_45_clk _00923_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__B _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload47 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10589_ net257 net2117 net423 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_8
Xclkload69 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload69/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__07957__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ top.lcd.cnt_500hz\[11\] _01449_ _06118_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12259_ _06080_ _06081_ net1119 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__o21a_1
XANTENNA__07148__B _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ top.DUT.register\[18\]\[31\] net778 net709 top.DUT.register\[7\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a22o_1
XANTENNA__13232__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06751_ top.DUT.register\[31\]\[28\] net803 net749 top.DUT.register\[1\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_75_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09470_ top.pc\[21\] _04494_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__nor2_1
X_06682_ _01778_ _01798_ net826 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_69_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08421_ net288 _03399_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or2_2
XANTENNA__06696__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ net905 top.pc\[3\] _03291_ _03465_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07303_ top.DUT.register\[17\]\[1\] net777 _02419_ vssd1 vssd1 vccd1 vccd1 _02420_
+ sky130_fd_sc_hd__a21o_1
X_08283_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload8 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload8/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout135_A _04208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ top.DUT.register\[13\]\[8\] net790 net717 top.DUT.register\[9\]\[8\] _02350_
+ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07165_ top.DUT.register\[26\]\[12\] net719 net580 top.DUT.register\[4\]\[12\] _02281_
+ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a221o_1
XANTENNA__10464__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_A _01856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1044_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07096_ top.DUT.register\[15\]\[15\] net806 net802 top.DUT.register\[31\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
XANTENNA__10952__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876__1136 vssd1 vssd1 vccd1 vccd1 _13876__1136/HI net1136 sky130_fd_sc_hd__conb_1
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 _04823_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout223 net225 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout671_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _04772_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 net247 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_208_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout256 _04753_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout769_A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 _04750_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
X_09806_ net208 top.DUT.register\[1\]\[14\] net390 vssd1 vssd1 vccd1 vccd1 _00136_
+ sky130_fd_sc_hd__mux2_1
Xfanout278 _01857_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout289 net291 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
X_07998_ top.DUT.register\[19\]\[21\] net672 _03112_ _03114_ vssd1 vssd1 vccd1 vccd1
+ _03115_ sky130_fd_sc_hd__a211o_1
XANTENNA__07581__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ net820 _04231_ net817 top.pc\[3\] vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a2bb2o_1
X_06949_ _02060_ _02061_ _02063_ _02065_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08125__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09668_ _04678_ _04686_ _04688_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or3_1
XANTENNA__07333__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ net396 _02639_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__nor2_1
XANTENNA__10639__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net353 _04607_ _04604_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__Y _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _05462_ _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__or2_1
XANTENNA__06418__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11561_ _05396_ _05416_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__xor2_4
XFILLER_0_80_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ clknet_leaf_99_clk _00846_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10512_ net169 net1702 net380 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _05284_ _05299_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13231_ clknet_leaf_22_clk _00777_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10374__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ net1541 net180 net510 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08061__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ clknet_leaf_2_clk _00708_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ net1489 net188 net430 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
X_12113_ _05971_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ clknet_leaf_47_clk _00639_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_12044_ _05853_ _05870_ _05856_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_53_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__B1 _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__X _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08116__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ clknet_leaf_106_clk _00492_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07324__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09864__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07712__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12877_ clknet_leaf_115_clk _00423_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10549__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ _05682_ _05686_ _05653_ _05668_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_190_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12848__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11759_ _05586_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload103 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_8
XFILLER_0_126_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ clknet_leaf_101_clk _00975_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06850__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _04013_ _04056_ _02928_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08689__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ top.DUT.register\[23\]\[25\] net567 net546 top.DUT.register\[24\]\[25\] _03037_
+ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a221o_1
XANTENNA_wire358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09552__A1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ top.DUT.register\[2\]\[26\] net685 net554 top.DUT.register\[22\]\[26\] _02968_
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a221o_1
XANTENNA__07563__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ _01919_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__inv_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_07783_ _02890_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__nor2_4
Xclkbuf_leaf_48_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08107__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _04551_ _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__and2b_1
X_06734_ top.DUT.register\[15\]\[3\] net689 net566 top.DUT.register\[23\]\[3\] _01850_
+ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07315__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06669__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _04472_ _04473_ _04471_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__o21ai_2
X_06665_ top.DUT.register\[13\]\[1\] net678 net670 top.DUT.register\[31\]\[1\] _01781_
+ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a221o_1
XANTENNA__10459__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08404_ net306 _03515_ _03500_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09384_ _04419_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_135_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06596_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__inv_2
XFILLER_0_191_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08335_ net315 _03448_ _03446_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout517_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08291__A1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ net394 _03357_ _03374_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a211o_2
XFILLER_0_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07094__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07217_ top.DUT.register\[14\]\[9\] net794 net586 top.DUT.register\[24\]\[9\] _02333_
+ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10194__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06841__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__B _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ _03311_ _03312_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09983__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09836__X _04833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ net322 _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_A _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A1 _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ net323 net351 _02176_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_144_Left_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09284__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ net246 net2172 net388 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 net1009 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07554__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12800_ clknet_leaf_14_clk _00346_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ clknet_leaf_64_clk _01305_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10992_ top.edg2.flip1 _01390_ _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and3_1
XFILLER_0_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07306__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12731_ clknet_leaf_1_clk _00277_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ clknet_leaf_104_clk _00208_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _05443_ net207 vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ clknet_leaf_7_clk _00139_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09459__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ _05387_ _05388_ net248 vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06832__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11475_ _05312_ _05315_ _05330_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or3b_1
XANTENNA__11169__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13214_ clknet_leaf_39_clk _00760_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ net1365 net255 net511 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_162_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13145_ clknet_leaf_42_clk _00691_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10832__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ net1379 net259 net431 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13076_ clknet_leaf_100_clk _00622_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10288_ net1595 net243 net522 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__mux2_1
X_12027_ _05849_ _05856_ _05864_ _05853_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_183_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06899__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_171_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ clknet_leaf_42_clk _00475_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10279__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13875__1135 vssd1 vssd1 vccd1 vccd1 _13875__1135/HI net1135 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_157_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06450_ net809 _01558_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__nor2_2
XFILLER_0_201_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06520__A1 top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06381_ top.d_ready _01493_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__or3_2
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ top.DUT.register\[30\]\[16\] net695 net679 top.DUT.register\[26\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a22o_1
XANTENNA__07076__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ top.DUT.register\[26\]\[23\] net679 net647 top.DUT.register\[12\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_180_Left_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07002_ top.DUT.register\[10\]\[19\] net726 net707 top.DUT.register\[7\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09773__A1 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06587__A1 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04020_ _04039_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_168_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09525__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ top.DUT.register\[1\]\[24\] net706 net562 top.DUT.register\[20\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ net473 _03970_ _03971_ net471 _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_90_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07000__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ net826 _02951_ _02617_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07766_ top.DUT.register\[30\]\[30\] net698 net563 top.DUT.register\[20\]\[30\] _02882_
+ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__a221o_1
XANTENNA__07352__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ top.pc\[23\] _04525_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11096__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__inv_2
XANTENNA__10189__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07697_ top.DUT.register\[4\]\[12\] net548 net623 top.DUT.register\[16\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09436_ _04470_ _04471_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_121_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06648_ top.DUT.register\[22\]\[2\] net553 net545 top.DUT.register\[24\]\[2\] _01764_
+ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09367_ _04405_ _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout801_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ _01676_ net799 _01662_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__and3b_4
XFILLER_0_170_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08318_ _03430_ _03431_ net288 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07067__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _02326_ _02775_ _04329_ _04330_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06814__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _01712_ _03281_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11260_ net901 _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ net169 net1799 net441 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
X_11191_ top.a1.halfData\[5\] net907 _01423_ _01427_ _01406_ vssd1 vssd1 vccd1 vccd1
+ _05098_ sky130_fd_sc_hd__o32a_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07775__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ net166 net1886 net444 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10073_ net170 top.DUT.register\[4\]\[23\] net446 vssd1 vssd1 vccd1 vccd1 _00241_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_42_clk _01355_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09461__B _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11087__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ clknet_leaf_73_clk _01288_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10099__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10975_ net1861 net165 net484 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12714_ clknet_leaf_116_clk _00260_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13694_ clknet_leaf_79_clk _00013_ net1088 vssd1 vssd1 vccd1 vccd1 top.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12645_ clknet_leaf_40_clk _00191_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10827__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12576_ clknet_leaf_15_clk _00122_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12327__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11527_ _05338_ _05384_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__xor2_2
XANTENNA__06805__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold309 top.DUT.register\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ _05287_ _05291_ _05296_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09755__A1 _03581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ net1431 net180 net514 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__mux2_1
XANTENNA__10562__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06612__Y _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11389_ _05228_ _05230_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07766__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ clknet_leaf_24_clk _00674_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13059_ clknet_leaf_34_clk _00605_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 top.DUT.register\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07518__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07620_ top.DUT.register\[26\]\[11\] net680 net668 top.DUT.register\[31\]\[11\] _02736_
+ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_163_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ top.a1.instruction\[30\] net857 _02667_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09140__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06502_ _01609_ _01618_ _01606_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_196_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07297__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ top.DUT.register\[23\]\[7\] net566 _02596_ _02598_ vssd1 vssd1 vccd1 vccd1
+ _02599_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _04268_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06433_ _01524_ _01542_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__nand2_1
XANTENNA__10737__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _04198_ _04202_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06364_ top.a1.instruction\[6\] _01486_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__nand2b_2
XANTENNA__06516__A top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08103_ top.DUT.register\[24\]\[22\] net545 net636 top.DUT.register\[25\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08797__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ net308 _03752_ _03772_ _03793_ _03727_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_79_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06295_ top.ramload\[21\] net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06235__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _03141_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or2_2
XANTENNA__09386__X _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08731__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold810 top.DUT.register\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 top.DUT.register\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 top.DUT.register\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold843 top.DUT.register\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10472__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 top.DUT.register\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 top.DUT.register\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold876 top.a1.row1\[60\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 top.DUT.register\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 top.DUT.register\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net251 net2294 net452 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout584_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _01878_ _02953_ _02957_ _04000_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07509__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09562__A _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ net1303 net861 net838 _03958_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout751_A _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09256__C_N _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ top.DUT.register\[17\]\[28\] net652 net632 top.DUT.register\[27\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a22o_1
X_08798_ _03129_ _03845_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07749_ top.DUT.register\[1\]\[31\] net706 net689 top.DUT.register\[15\]\[31\] _02865_
+ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07288__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ net235 net2080 net372 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07810__A _01898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ top.pc\[18\] _04445_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or2_1
X_10691_ top.DUT.register\[23\]\[5\] net251 net500 vssd1 vssd1 vccd1 vccd1 _00831_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10647__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12430_ clknet_leaf_78_clk top.ru.next_FetchedData\[25\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12361_ net2166 _06141_ net814 vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07996__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ net901 _05165_ _05178_ _05180_ net845 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12292_ net1782 _06100_ net1118 vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06713__X _01830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07460__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11243_ net871 _05039_ _05049_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and3_1
XANTENNA__10382__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13874__1134 vssd1 vssd1 vccd1 vccd1 _13874__1134/HI net1134 sky130_fd_sc_hd__conb_1
XANTENNA__06161__A top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07212__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net63 net885 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__and2_1
X_10125_ net239 net2096 net445 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10056_ net244 top.DUT.register\[4\]\[6\] net448 vssd1 vssd1 vccd1 vccd1 _00224_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08173__B1 _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08088__A _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ clknet_leaf_72_clk _01340_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13746_ clknet_leaf_67_clk _01271_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07279__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ net1514 net235 net483 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10557__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13677_ clknet_leaf_75_clk _01218_ net1082 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
X_10889_ net2206 net249 net408 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ clknet_leaf_98_clk _00174_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08779__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ clknet_leaf_86_clk _00105_ net1019 vssd1 vssd1 vccd1 vccd1 top.pc\[24\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 top.DUT.register\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07451__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold117 top.ramstore\[18\] vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top.pad.button_control.r_counter\[14\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10292__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
XANTENNA__08400__B2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 _04343_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _03623_ net456 net535 _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__o211a_2
X_06982_ _02092_ _02094_ _02096_ _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__or4_4
XANTENNA_wire340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ net461 _03803_ _03808_ net466 _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A1 top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ net394 _03744_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__nand2_1
XANTENNA__06714__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ _02718_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__nand2_2
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08583_ net472 _03684_ _03687_ _02522_ _03678_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_A _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07534_ top.DUT.register\[17\]\[13\] net651 net639 top.DUT.register\[9\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08285__X _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10467__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07465_ top.DUT.register\[13\]\[6\] net677 net641 top.DUT.register\[9\]\[6\] _02581_
+ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1074_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09204_ top.pc\[5\] _04239_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__and2_1
X_06416_ net810 _01532_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07396_ net285 _02409_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07690__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ _01612_ _04185_ _04186_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__and4_1
X_06347_ _01332_ _01468_ _01333_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07978__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _03407_ _04118_ _03441_ _03516_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__or4b_1
XFILLER_0_32_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06278_ net1221 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[4\] sky130_fd_sc_hd__and2_1
XANTENNA__08461__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ top.DUT.register\[15\]\[19\] net687 net675 top.DUT.register\[13\]\[19\] _03133_
+ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a221o_1
XANTENNA__06650__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 top.DUT.register\[17\]\[27\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 top.DUT.register\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08180__B _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold662 top.DUT.register\[17\]\[29\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 top.DUT.register\[9\]\[10\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _01183_ vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 top.DUT.register\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _04944_ _04945_ _04942_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__o21ai_1
X_08919_ net274 _03472_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nor2_1
XANTENNA__12714__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ _04557_ net360 net328 top.a1.dataIn\[24\] net363 vssd1 vssd1 vccd1 vccd1
+ _04889_ sky130_fd_sc_hd__a221o_1
X_11930_ _05714_ _05752_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nor2_1
XANTENNA__07902__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11861_ _05720_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__nor2_1
X_13600_ clknet_leaf_55_clk _01141_ net1095 vssd1 vssd1 vccd1 vccd1 top.ramload\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10812_ net155 net1282 net410 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08458__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ _05618_ _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ clknet_leaf_0_clk _01077_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10743_ net167 net2274 net417 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10377__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06427__Y _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13462_ clknet_leaf_105_clk _01008_ net981 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10674_ net179 net1893 net419 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12413_ clknet_leaf_54_clk top.ru.next_FetchedData\[8\] net1099 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[8\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_209_Right_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13502__RESET_B net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13393_ clknet_leaf_8_clk _00939_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07969__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ _01506_ _01507_ _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06443__X _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06641__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12275_ top.lcd.cnt_20ms\[8\] _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__and2_1
X_11226_ _01418_ net405 _04682_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10840__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net923 net1304 net875 _05078_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ net167 net2174 net389 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output59_A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ net1219 net883 net848 top.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a22o_1
XANTENNA__09343__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ net163 net2093 net531 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
XANTENNA__07434__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06618__X _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07450__A _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ clknet_leaf_63_clk _01259_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ net321 _02366_ _02347_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06201_ net908 net909 top.a1.state\[0\] vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__or3b_1
XANTENNA__06880__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ _02291_ _02293_ _02295_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07424__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08281__A _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout405 _05107_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_2
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_6
XFILLER_0_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout427 net429 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
X_09822_ _04199_ _04763_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nor2_1
XANTENNA__10750__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _04976_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_6
Xfanout449 _04967_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07625__A _02305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ net820 _04279_ top.a1.dataIn\[7\] net813 vssd1 vssd1 vccd1 vccd1 _04760_
+ sky130_fd_sc_hd__a2bb2o_1
X_06965_ top.DUT.register\[3\]\[21\] net782 net775 top.DUT.register\[2\]\[21\] _02081_
+ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _03106_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__xnor2_2
X_09684_ _04701_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nor2_1
X_06896_ _02006_ _02008_ _02010_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or4_2
XFILLER_0_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09796__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08635_ net463 _03718_ _03731_ _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_87_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06699__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout547_A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07631__Y _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ _02743_ _03648_ _02744_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a21boi_1
XANTENNA__08456__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07517_ top.DUT.register\[6\]\[14\] net576 net671 top.DUT.register\[19\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
XANTENNA__10197__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ _02772_ _03584_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__nand2_1
X_13873__1133 vssd1 vssd1 vccd1 vccd1 _13873__1133/HI net1133 sky130_fd_sc_hd__conb_1
XANTENNA_fanout714_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09986__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07448_ _02526_ _02564_ net401 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
XANTENNA__07663__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06871__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ top.DUT.register\[5\]\[4\] net602 net768 top.DUT.register\[11\]\[4\] _02495_
+ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10925__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13654__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ net857 _01632_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__or2_4
XANTENNA__07415__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net1603 net258 net514 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__mux2_1
XANTENNA__08612__B2 _03715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09049_ _04065_ _04101_ _03960_ _04045_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__and4b_1
XANTENNA__07078__Y _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__12966__RESET_B net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06423__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ _05919_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__nand2_1
Xhold470 top.DUT.register\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 top.DUT.register\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 _01186_ vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net1170 _05028_ net480 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
XANTENNA__10660__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net960 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_2
Xfanout961 net969 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 net978 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08128__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09325__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout994 net1021 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_11_clk _00508_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1170 top.pad.keyCode\[6\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net125 net126 _05744_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a21oi_2
Xhold1181 top.DUT.register\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11683__B1 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1192 top.DUT.register\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ clknet_leaf_120_clk _00439_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_206_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11844_ _05660_ _05694_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12227__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06438__X _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ _05612_ _05614_ _05594_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09896__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10726_ net237 net2064 net416 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
X_13514_ clknet_leaf_117_clk _01060_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13445_ clknet_leaf_40_clk _00991_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06862__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10835__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ net255 net1466 net421 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09909__B _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload15 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__09197__A _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload26 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08603__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload37 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_8
X_13376_ clknet_leaf_13_clk _00922_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10588_ net262 net1928 net424 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload48 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__clkinv_8
Xclkload59 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload59/X sky130_fd_sc_hd__clkbuf_4
X_12327_ _06122_ net742 _06121_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12258_ top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _06081_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11209_ _05018_ _05033_ net369 net404 net1267 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a32o_1
XANTENNA__10570__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ _06043_ _06044_ _06048_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__or3_1
XFILLER_0_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06917__A1 top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06750_ top.DUT.register\[13\]\[28\] net789 net585 top.DUT.register\[24\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06681_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ net281 _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07893__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08351_ net395 _03441_ _03464_ net470 _03458_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__a221o_4
XFILLER_0_129_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07302_ top.DUT.register\[15\]\[1\] net807 net803 top.DUT.register\[31\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22o_1
XANTENNA__13677__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08282_ net318 _01984_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08563__X _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07645__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XFILLER_0_74_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06853__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07233_ top.DUT.register\[14\]\[8\] net794 net709 top.DUT.register\[7\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a22o_1
XANTENNA__10745__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__A1 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ top.DUT.register\[31\]\[12\] net800 net770 top.DUT.register\[27\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08070__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07095_ _02205_ _02207_ _02209_ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout202 _04823_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_1
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 net215 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_1
Xfanout235 _04772_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_1
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _03738_ net454 net533 _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o211a_1
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
Xfanout268 _04750_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_1
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
X_07997_ top.DUT.register\[7\]\[21\] net574 net570 top.DUT.register\[21\]\[21\] _03113_
+ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06948_ top.DUT.register\[24\]\[22\] net585 net712 top.DUT.register\[25\]\[22\] _02064_
+ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a221o_1
X_09736_ net258 net1570 net390 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09667_ top.a1.state\[0\] _04687_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _00113_
+ sky130_fd_sc_hd__o22a_1
X_06879_ top.DUT.register\[1\]\[25\] net780 net717 top.DUT.register\[9\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout831_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08618_ _03617_ _03719_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09598_ _04623_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08549_ net303 _03654_ _03653_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06418__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _05394_ _05411_ _05412_ _05392_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07636__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ net173 net1672 net378 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
XANTENNA__10655__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _05342_ _05345_ _05348_ _05349_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230_ clknet_leaf_94_clk _00776_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10442_ net1448 net183 net510 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13161_ clknet_leaf_27_clk _00707_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08061__A2 _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10373_ net1442 net193 net430 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
X_12112_ _05958_ _05964_ _05959_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13092_ clknet_leaf_29_clk _00638_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12043_ _05892_ _05894_ _05869_ _05871_ _05883_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10390__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07572__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
Xfanout791 _01530_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07552__X _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09480__A _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_10_clk _00491_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08521__B1 _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07712__B _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12876_ clknet_leaf_115_clk _00422_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11827_ _05682_ _05686_ _05668_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_190_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07088__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ _05612_ _05614_ _05590_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ net1660 net173 net498 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XANTENNA__06835__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10565__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12888__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11689_ _05518_ _05536_ _05539_ _05529_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_155_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload104 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_155_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13428_ clknet_leaf_99_clk _00974_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13359_ clknet_leaf_20_clk _00905_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08052__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07260__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ top.DUT.register\[17\]\[25\] net654 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__and2_1
XANTENNA__09001__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872__1132 vssd1 vssd1 vccd1 vccd1 _13872__1132/HI net1132 sky130_fd_sc_hd__conb_1
X_07851_ top.DUT.register\[30\]\[26\] net697 net550 top.DUT.register\[4\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06802_ _01909_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__nor2_8
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_1
X_07782_ _02892_ _02894_ _02896_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__or4_2
XFILLER_0_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ top.pc\[24\] _02615_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or2_1
X_06733_ top.DUT.register\[19\]\[3\] net673 net653 top.DUT.register\[17\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
XANTENNA__13605__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__inv_2
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06664_ top.DUT.register\[30\]\[1\] net698 net686 top.DUT.register\[2\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08403_ net301 _03514_ _03502_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a21o_1
XANTENNA__09068__A1 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ _04420_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__and2b_1
X_06595_ net366 net326 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ _03447_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07618__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08265_ _03326_ _03380_ net471 vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10475__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout412_A _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ top.DUT.register\[9\]\[9\] net717 net759 top.DUT.register\[2\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ net300 net334 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__and2_1
XANTENNA__12558__RESET_B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07147_ net365 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__inv_2
XANTENNA__08043__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__Y _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07078_ net350 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__inv_2
XANTENNA__09791__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout879_A _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09284__B _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1019 net1020 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XANTENNA__07003__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07085__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13842__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09719_ _04729_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_1
X_10991_ _05005_ _05007_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ clknet_leaf_20_clk _00276_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07857__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12661_ clknet_leaf_101_clk _00207_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _05470_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_172_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ clknet_leaf_116_clk _00138_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07609__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11543_ top.a1.dataIn\[14\] _05401_ _05402_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10385__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12981__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07490__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11474_ _05313_ _05330_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ clknet_leaf_119_clk _00759_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ net1330 net266 net511 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13144_ clknet_leaf_33_clk _00690_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ net1534 net261 net432 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_108_clk _00621_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ _04183_ net615 _04973_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_4
XANTENNA__06611__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_183_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07723__A _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12928_ clknet_leaf_13_clk _00474_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07848__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_1_clk _00405_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06380_ _01499_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06808__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08050_ top.DUT.register\[25\]\[23\] net635 _03164_ _03166_ vssd1 vssd1 vccd1 vccd1
+ _03167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07481__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07001_ top.DUT.register\[21\]\[19\] net608 net596 top.DUT.register\[6\]\[19\] _02117_
+ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08025__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07233__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07784__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__B1 _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ _04020_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_168_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ top.DUT.register\[8\]\[24\] net559 net666 top.DUT.register\[14\]\[24\] _03019_
+ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08883_ net279 _02518_ _03403_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_205_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ _02941_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__or2_2
XFILLER_0_169_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07765_ top.DUT.register\[26\]\[30\] net682 net678 top.DUT.register\[13\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a22o_1
XANTENNA__09289__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08448__B _01856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11096__A1 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ top.pc\[23\] _04525_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nor2_1
X_06716_ top.a1.instruction\[24\] net855 _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__o21a_1
X_07696_ top.DUT.register\[23\]\[12\] net564 net640 top.DUT.register\[9\]\[12\] _02812_
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a221o_1
XANTENNA__06249__A top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09435_ top.pc\[19\] _04460_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__nand2_1
X_06647_ top.DUT.register\[12\]\[2\] net649 net628 top.DUT.register\[29\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _04385_ _04386_ _04387_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__o21ai_2
X_06578_ net747 _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ _03308_ _03320_ net320 vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09279__B _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _04339_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08183__B _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09994__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ net465 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08016__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ net1337 net860 _03294_ net837 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
X_10210_ net170 net2108 net438 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07224__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net1376 _05097_ _05096_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
XANTENNA__06712__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net171 net1817 net442 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XANTENNA__09516__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ net177 net2335 net447 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XANTENNA__08724__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ clknet_leaf_42_clk net1251 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09461__C _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06750__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ clknet_leaf_66_clk _01287_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ net1655 net166 net483 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ clknet_leaf_27_clk _00259_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13693_ clknet_leaf_79_clk _00007_ net1087 vssd1 vssd1 vccd1 vccd1 top.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_183_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06593__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ clknet_leaf_28_clk _00190_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13871__1131 vssd1 vssd1 vccd1 vccd1 _13871__1131/HI net1131 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_61_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ clknet_leaf_77_clk _00121_ net1080 vssd1 vssd1 vccd1 vccd1 top.pc\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07463__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11526_ top.a1.dataIn\[15\] _05384_ _05385_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__or3_1
XANTENNA__08661__X _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10843__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08007__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _05287_ _05296_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__nand2_2
XFILLER_0_150_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10408_ net2152 net186 net514 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__mux2_1
XANTENNA__07215__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07718__A _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06622__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11388_ _05221_ _05225_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10339_ net1589 net196 net518 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
X_13127_ clknet_leaf_49_clk _00673_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13058_ clknet_leaf_10_clk _00604_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12009_ _05849_ _05864_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ _01641_ _01777_ net401 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_200_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09140__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06501_ _01487_ _01611_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__o21ai_1
X_07481_ top.DUT.register\[5\]\[7\] net542 net653 top.DUT.register\[17\]\[7\] _02597_
+ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _01412_ _02528_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__xnor2_1
X_06432_ net812 _01532_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_17_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _04079_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06363_ _01483_ net914 top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ top.DUT.register\[30\]\[22\] net696 net541 top.DUT.register\[5\]\[22\] _03218_
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07454__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ _03854_ _03873_ _03888_ _03910_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_79_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08797__A3 _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06294_ net1297 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[20\] sky130_fd_sc_hd__and2_1
XFILLER_0_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08033_ _03143_ _03145_ _03147_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__or4_1
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10753__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold800 top.DUT.register\[9\]\[8\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 top.DUT.register\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout208_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__Y _01920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold822 top.DUT.register\[29\]\[26\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09746__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 top.DUT.register\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 top.DUT.register\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold855 top.DUT.register\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 top.DUT.register\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 top.DUT.register\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 top.DUT.register\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 top.DUT.register\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net253 net2327 net452 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__mux2_1
XANTENNA__06251__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ net1294 net860 net837 _04023_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__a22o_1
XANTENNA__06980__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09562__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ top.ru.state\[5\] top.pc\[25\] net539 _03957_ vssd1 vssd1 vccd1 vccd1 _03958_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08459__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07817_ top.DUT.register\[7\]\[28\] net574 net685 top.DUT.register\[2\]\[28\] _02933_
+ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a221o_1
X_08797_ net310 net470 _03541_ _03889_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__a311o_1
XFILLER_0_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06732__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ top.DUT.register\[17\]\[31\] net653 net633 top.DUT.register\[27\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ _02776_ _02795_ net825 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10928__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout911_A top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08906__B _03995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07810__B _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ top.pc\[18\] _04445_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07693__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ net2188 net253 net499 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_3__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ net841 _01748_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12360_ top.pad.button_control.r_counter\[6\] _06141_ vssd1 vssd1 vccd1 vccd1 _06143_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_43_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11311_ top.a1.row1\[122\] _05129_ _05138_ top.a1.row2\[10\] _05179_ vssd1 vssd1
+ vccd1 vccd1 _05180_ sky130_fd_sc_hd__a221o_1
XANTENNA__06799__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ top.lcd.cnt_20ms\[14\] _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2_1
XANTENNA__10663__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__Y _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ _05121_ net1231 net403 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ net924 net1301 net876 _05086_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ net244 net1683 net444 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ net250 net1920 net448 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06723__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ clknet_leaf_72_clk _01339_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_11_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08656__X _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13745_ clknet_leaf_67_clk _01270_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10838__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ net1795 net237 net484 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07684__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08308__S _01856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ clknet_leaf_88_clk _01217_ net1082 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
X_10888_ net1684 net256 net408 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ clknet_leaf_111_clk _00173_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12558_ clknet_leaf_85_clk _00104_ net1019 vssd1 vssd1 vccd1 vccd1 top.pc\[23\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08832__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10573__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ _05299_ _05332_ _05298_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 top.a1.row1\[19\] vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ clknet_leaf_90_clk _00036_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold118 top.a1.row1\[112\] vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 top.ramaddr\[26\] vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12504__D net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__A2 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net611 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ top.DUT.register\[22\]\[20\] net605 net776 top.DUT.register\[17\]\[20\] _02097_
+ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_14__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _03816_ _03817_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__and3_1
XANTENNA__09382__B _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08651_ net474 net309 _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_198_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A2 _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06714__A2 _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _02222_ _02715_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net309 _03686_ _03673_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07470__X _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07533_ top.DUT.register\[25\]\[13\] net635 _02647_ _02649_ vssd1 vssd1 vccd1 vccd1
+ _02650_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10748__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout158_A _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07675__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ top.DUT.register\[26\]\[6\] net681 net658 top.DUT.register\[28\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ net918 top.pc\[4\] _04253_ top.testpc.en_latched vssd1 vssd1 vccd1 vccd1
+ _00085_ sky130_fd_sc_hd__o211a_1
X_06415_ _01520_ _01527_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07395_ _01737_ net285 _02429_ net289 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06246__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ top.a1.instruction\[28\] top.a1.instruction\[29\] top.a1.instruction\[30\]
+ top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__and4_1
X_06346_ _01332_ _01472_ _01476_ _01462_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XANTENNA__07427__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ net310 _03686_ _03903_ _03929_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__a2111o_1
X_06277_ net1902 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[3\] sky130_fd_sc_hd__and2_1
XANTENNA__10483__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08461__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ top.DUT.register\[17\]\[19\] net651 net623 top.DUT.register\[16\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold630 top.DUT.register\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 top.DUT.register\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 top.DUT.register\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 top.DUT.register\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold674 top.DUT.register\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 top.DUT.register\[28\]\[17\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 top.DUT.register\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ net144 top.DUT.register\[1\]\[30\] net393 vssd1 vssd1 vccd1 vccd1 _00152_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout861_A _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net308 _03683_ _03852_ net271 _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__o221a_1
X_13870__1130 vssd1 vssd1 vccd1 vccd1 _13870__1130/HI net1130 sky130_fd_sc_hd__conb_1
XANTENNA__08155__A1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net820 _04548_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_1
X_08849_ _03327_ _03346_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06705__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _05677_ _05709_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ net158 net2091 net411 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__mux2_1
XANTENNA__10658__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ _05629_ _05630_ net129 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_45_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07666__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ clknet_leaf_16_clk _01076_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10742_ net171 net2169 net414 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06437__A top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07130__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ net183 net1925 net418 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__mux2_1
X_13461_ clknet_leaf_101_clk _01007_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07418__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ clknet_leaf_54_clk top.ru.next_FetchedData\[7\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08652__A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ clknet_leaf_117_clk _00938_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12343_ top.pad.button_control.debounce top.pad.button_control.noisy vssd1 vssd1
+ vccd1 vccd1 _06132_ sky130_fd_sc_hd__nand2_1
XANTENNA__10393__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ _06090_ net1117 _06089_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11225_ net1254 net404 net369 _05113_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a22o_1
XANTENNA__10725__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ net53 net880 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06944__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ net172 net1774 net386 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ net100 net886 net849 net1234 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__a22o_1
XANTENNA__09770__X _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ net167 net2083 net531 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XANTENNA__12410__Q top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09930__B _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10568__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _05831_ _05842_ _05843_ _05847_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__or4b_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ clknet_leaf_62_clk _01258_ net1109 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[15\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_193_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13659_ clknet_leaf_89_clk _01200_ net1015 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
X_06200_ top.a1.state\[2\] net909 top.a1.state\[0\] vssd1 vssd1 vccd1 vccd1 _01420_
+ sky130_fd_sc_hd__nor3b_2
XFILLER_0_128_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07180_ top.DUT.register\[5\]\[11\] net601 net716 top.DUT.register\[9\]\[11\] _02296_
+ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08082__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__Y _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06632__B2 top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08909__B1 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net409 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout417 _04996_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12480__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ net818 _04433_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__nor2_1
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_6
Xfanout439 _04976_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_4
XANTENNA__06935__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ net245 net1547 net392 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
X_06964_ top.DUT.register\[18\]\[21\] net779 net767 top.DUT.register\[11\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08703_ _03207_ _03784_ _03206_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__o21a_1
X_09683_ top.pad.keyCode\[5\] top.pad.keyCode\[6\] top.pad.keyCode\[7\] top.pad.keyCode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__or4b_2
X_06895_ top.DUT.register\[28\]\[24\] net741 net582 top.DUT.register\[4\]\[24\] _02011_
+ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a221o_1
XANTENNA__09885__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07896__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ net467 _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__B _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07360__A2 _01545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ net1421 net858 net836 _03670_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09637__A1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07516_ top.DUT.register\[4\]\[14\] net548 net655 top.DUT.register\[28\]\[14\] _02632_
+ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__a221o_1
XANTENNA__07648__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ net1306 net860 net837 _03604_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07112__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ top.a1.instruction\[19\] _01616_ _01640_ top.a1.instruction\[27\] vssd1 vssd1
+ vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_2
XFILLER_0_146_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06320__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07378_ top.DUT.register\[25\]\[4\] net713 net709 top.DUT.register\[7\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06329_ _01459_ _01332_ _01331_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__mux2_1
X_09117_ net856 _01632_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nor2_2
XANTENNA__08073__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__A2 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__B _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ _03982_ _04001_ _04025_ _04100_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__and4_1
XANTENNA__07820__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 top.DUT.register\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 top.DUT.register\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ top.a1.dataIn\[3\] net869 _05005_ _05027_ vssd1 vssd1 vccd1 vccd1 _05028_
+ sky130_fd_sc_hd__a211o_1
Xhold482 top.DUT.register\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 top.DUT.register\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06926__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net942 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
Xfanout951 net959 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
Xfanout962 net969 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12935__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout973 net978 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_2
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout995 net998 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ clknet_leaf_45_clk _00507_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1160 top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1171 top.DUT.register\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _05768_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__and2_1
Xhold1182 top.DUT.register\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07887__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 top.DUT.register\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ clknet_leaf_51_clk _00438_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_206_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _05666_ _05691_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10388__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07639__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ _05593_ _05617_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__xor2_2
XANTENNA__07103__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ clknet_leaf_27_clk _01059_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10725_ net245 net1736 net416 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09478__A _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13444_ clknet_leaf_29_clk _00990_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ net267 net1439 net421 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_6
XANTENNA__09197__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13375_ clknet_leaf_32_clk _00921_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10587_ net241 net1954 net423 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__mux2_1
Xclkload27 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload38 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__06614__B net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload49 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_8
XFILLER_0_152_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[10\] _06118_ vssd1 vssd1 vccd1
+ vccd1 _06122_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12405__Q top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ _01384_ _06080_ net1119 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o21a_1
XANTENNA__10851__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08367__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _05015_ _05029_ net369 net405 net1249 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a32o_1
XANTENNA__07726__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12188_ _06044_ _06048_ _06043_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06917__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ net922 net1536 net874 _05069_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07590__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06680_ _01787_ _01796_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__or2_4
XANTENNA__07878__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06629__X _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10298__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08844__X _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07301_ _02411_ _02413_ _02415_ _02417_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__or4_2
XFILLER_0_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ _01800_ _01879_ _01899_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08842__A2 _03927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07232_ top.DUT.register\[22\]\[8\] net606 net774 top.DUT.register\[2\]\[8\] _02348_
+ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08055__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ top.DUT.register\[12\]\[12\] net734 _02278_ _02279_ vssd1 vssd1 vccd1 vccd1
+ _02280_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07802__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ top.DUT.register\[5\]\[15\] net602 net764 top.DUT.register\[19\]\[15\] _02210_
+ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10761__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout203 _04814_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
Xfanout225 net227 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _04762_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
X_09804_ net816 _04803_ _04797_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a21o_1
Xfanout247 _04759_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ top.DUT.register\[3\]\[21\] net692 net676 top.DUT.register\[13\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__a22o_1
XANTENNA__07581__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _03425_ net456 net535 _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__o211a_2
X_06947_ top.DUT.register\[27\]\[22\] net771 net589 top.DUT.register\[20\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _04675_ net872 _04684_ _04686_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a211o_1
X_06878_ top.DUT.register\[22\]\[25\] net606 _01994_ vssd1 vssd1 vccd1 vccd1 _01995_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07333__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ _03533_ _03570_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _04622_ _01878_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__and2b_1
XFILLER_0_139_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09997__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ net283 _03461_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10936__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ net282 _02028_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10510_ net176 net1735 net379 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
XANTENNA__09025__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11490_ _05346_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ net1345 net188 net510 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08046__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09794__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ net1978 net197 net431 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
X_13160_ clknet_leaf_24_clk _00706_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12111_ _05960_ _05963_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13091_ clknet_leaf_34_clk _00637_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10671__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12042_ _05892_ _05894_ _05869_ _05883_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__a211o_1
XANTENNA__07546__A _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 top.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
Xfanout781 _01539_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
XANTENNA__09761__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout792 _01529_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09480__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ clknet_leaf_117_clk _00490_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ clknet_leaf_6_clk _00421_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11826_ _05682_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11757_ _05584_ _05616_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10846__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ net1434 net174 net497 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
XANTENNA__08316__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11688_ _05547_ _05548_ _05543_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06625__A _01733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload105 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__clkinv_2
X_13427_ clknet_leaf_110_clk _00973_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ net187 top.DUT.register\[21\]\[19\] net374 vssd1 vssd1 vccd1 vccd1 _00781_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__B1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_93_clk _00904_ net997 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12309_ top.lcd.cnt_500hz\[4\] _01447_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__or2_1
XANTENNA__10581__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13289_ clknet_leaf_9_clk _00835_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06360__A top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07850_ _02960_ _02962_ _02964_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__or4_1
XANTENNA__07563__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _01911_ _01913_ _01915_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_3_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07781_ top.DUT.register\[24\]\[30\] net547 net626 top.DUT.register\[16\]\[30\] _02897_
+ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a221o_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06771__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ top.pc\[24\] _02615_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__and2_1
XANTENNA__13644__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06732_ top.DUT.register\[20\]\[3\] net562 net547 top.DUT.register\[24\]\[3\] _01848_
+ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07315__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__B2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06663_ top.DUT.register\[3\]\[1\] net693 net662 top.DUT.register\[18\]\[1\] _01779_
+ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a221o_1
X_09451_ _04484_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08402_ _03401_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__or2_1
X_06594_ net323 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ _01415_ _04411_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09068__A2 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ net297 net340 _03311_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10756__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout238_A _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ net308 _03379_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nor2_1
XANTENNA__06826__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06535__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08028__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07215_ top.DUT.register\[18\]\[9\] net778 net724 top.DUT.register\[16\]\[9\] _02331_
+ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a221o_1
X_08195_ net322 net343 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__and2_1
XANTENNA__09225__C1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _02255_ _02258_ _02260_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__nor4_1
XANTENNA__09776__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10491__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07077_ _02187_ _02190_ _02191_ _02193_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__nor4_1
XFILLER_0_140_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12527__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1021 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA_fanout774_A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08200__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ top.DUT.register\[22\]\[18\] net552 net544 top.DUT.register\[24\]\[18\] _03095_
+ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07372__Y _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ top.a1.instruction\[8\] _04730_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__or2_1
XANTENNA__07813__B _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ net920 _05006_ net797 net865 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__o211a_1
XANTENNA__07306__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ _01417_ net853 _04224_ _04672_ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13386__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ clknet_leaf_99_clk _00206_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ _05439_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__xor2_1
XANTENNA__13315__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12591_ clknet_leaf_25_clk _00137_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_67_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _01395_ net248 _05386_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_208_Left_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08019__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09216__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ _05302_ _05331_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_137_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ clknet_leaf_16_clk _00758_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11169__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ net2036 net257 net509 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11574__B1 top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ clknet_leaf_114_clk _00689_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ net1690 net241 net431 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ net140 net2291 net437 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__mux2_1
X_13074_ clknet_leaf_104_clk _00620_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12025_ _05841_ _05865_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13667__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06753__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11526__A top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B _02549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09298__A2 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12927_ clknet_leaf_23_clk _00473_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12858_ clknet_leaf_15_clk _00404_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08835__A _02519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _05631_ net129 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_107_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ clknet_leaf_81_clk _00335_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ top.DUT.register\[26\]\[19\] net719 net580 top.DUT.register\[4\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07784__A2 _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ _04033_ _04035_ _04038_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_168_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07902_ top.DUT.register\[17\]\[24\] net653 net633 top.DUT.register\[27\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08882_ _02983_ _03371_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07914__A _02023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _02943_ _02945_ _02947_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__or4_1
XANTENNA__06744__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__Y _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_108_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09503_ top.pc\[23\] _04529_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__nor2_1
X_06715_ _01630_ _01750_ _01806_ net401 net856 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a221o_1
XANTENNA__11096__A2 _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ top.DUT.register\[19\]\[12\] net671 net652 top.DUT.register\[17\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06249__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ top.pc\[19\] _04460_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__nor2_1
X_06646_ _01756_ _01758_ _01760_ _01762_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09365_ _04403_ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10486__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ top.DUT.register\[24\]\[0\] net545 net660 top.DUT.register\[18\]\[0\] _01693_
+ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_191_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08316_ _03313_ _03323_ net285 vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09296_ _04323_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _01728_ _01736_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or2_1
XANTENNA__07472__A1 top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09749__B1 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ net905 top.ru.state\[0\] _01511_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout989_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ top.DUT.register\[15\]\[13\] net805 net800 top.DUT.register\[31\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06712__B _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ net174 net1763 net443 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XANTENNA__08972__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net182 net2046 net448 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__B1 _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_42_clk _01353_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11087__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ clknet_leaf_65_clk _01286_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10973_ net1623 net172 net482 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ clknet_leaf_26_clk _00258_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ clknet_leaf_79_clk _00012_ net1088 vssd1 vssd1 vccd1 vccd1 top.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12643_ clknet_leaf_35_clk _00189_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10396__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08374__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12574_ clknet_leaf_60_clk _00120_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[5\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_61_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06175__A top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ _05384_ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08390__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _05313_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__and2_1
X_10407_ net1521 net188 net513 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07718__B _02587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11387_ _05246_ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_185_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06622__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ clknet_leaf_22_clk _00672_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ net1739 net199 net517 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06974__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__Q top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__Y _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ clknet_leaf_49_clk _00603_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net209 net1707 net434 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07518__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _05848_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__xor2_2
XANTENNA__11256__A top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13237__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06500_ _01515_ net824 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__or2_1
X_07480_ top.DUT.register\[15\]\[7\] net689 net625 top.DUT.register\[16\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
XANTENNA__07151__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06637__X _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06431_ net809 _01543_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__nor2_4
XFILLER_0_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06362_ top.a1.instruction\[6\] _01483_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__or2_2
XFILLER_0_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ _04202_ _04198_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ top.DUT.register\[13\]\[22\] net676 net628 top.DUT.register\[29\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09081_ _03842_ _04115_ _04123_ _04128_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__o32a_1
X_06293_ net2307 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[19\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13832__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ top.DUT.register\[8\]\[19\] net556 net663 top.DUT.register\[14\]\[19\] _03148_
+ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold801 top.DUT.register\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 top.DUT.register\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 top.DUT.register\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold834 top.DUT.register\[26\]\[0\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold845 top.DUT.register\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold856 top.DUT.register\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 top.DUT.register\[28\]\[10\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 top.DUT.register\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ net267 net2243 net453 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__mux2_1
Xhold889 top.DUT.register\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ net904 top.pc\[28\] net538 _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a22o_1
XANTENNA__07509__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08865_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout472_A _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__B net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ top.DUT.register\[15\]\[28\] net690 net681 top.DUT.register\[26\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a22o_1
X_08796_ _01741_ _03230_ _03232_ net459 _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07390__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07747_ top.DUT.register\[14\]\[31\] net666 net550 top.DUT.register\[4\]\[31\] _02863_
+ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07650__Y _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07142__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _02785_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__nor2_2
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09417_ _04440_ _04441_ _04439_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21ai_2
X_06629_ _01719_ _01744_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__or2_2
XANTENNA__08890__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09348_ _04385_ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_101_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ top.pc\[10\] _02668_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__and2b_1
X_11310_ top.a1.row2\[2\] _05132_ _05134_ top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1
+ _05179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07996__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ _06100_ net1118 _06099_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_134_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12542__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ net872 _05035_ _05046_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07748__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ net61 net884 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and2_1
XANTENNA__06956__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ net250 net1948 net444 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ net255 net1444 net448 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06708__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A2 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07381__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_72_clk _01338_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13330__RESET_B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10268__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13744_ clknet_leaf_67_clk _01269_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10956_ net2121 net246 net483 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XANTENNA__07133__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13675_ clknet_leaf_90_clk _01216_ net1010 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
X_10887_ top.DUT.register\[29\]\[3\] net268 net408 vssd1 vssd1 vccd1 vccd1 _01021_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ clknet_leaf_106_clk _00172_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__X _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_159_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12408__Q top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10854__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12557_ clknet_leaf_85_clk _00103_ net1019 vssd1 vssd1 vccd1 vccd1 top.pc\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09928__B _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__B _03924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07729__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _05333_ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nor2_1
XANTENNA__08324__S _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ clknet_leaf_90_clk _00035_ net1011 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold108 net115 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 top.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ net327 _05295_ _05274_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06947__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13109_ clknet_leaf_101_clk _00655_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06980_ top.DUT.register\[6\]\[20\] net597 net581 top.DUT.register\[4\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13418__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08650_ _03565_ _03751_ net283 vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_198_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07601_ _02222_ _02715_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ _03674_ _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07532_ top.DUT.register\[22\]\[13\] net552 net647 top.DUT.register\[12\]\[13\] _02648_
+ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a221o_1
XANTENNA__07124__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ top.DUT.register\[23\]\[6\] net566 net685 top.DUT.register\[2\]\[6\] _02579_
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06527__B _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ net133 _04241_ _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06414_ net812 _01525_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__nor2_1
X_07394_ net289 _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ top.a1.instruction\[6\] top.a1.instruction\[20\] top.a1.instruction\[19\]
+ top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__and4_1
X_06345_ _01465_ _01472_ _01335_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10764__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout220_A _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07978__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06276_ net1947 net899 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[2\] sky130_fd_sc_hd__and2_1
X_09064_ net276 _03533_ _02518_ net356 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_115_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08234__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08015_ _03128_ _03129_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__and2b_2
XANTENNA__06650__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold620 top.ramload\[1\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 top.DUT.register\[27\]\[7\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06262__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap350 net352 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
Xhold642 top.DUT.register\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 top.DUT.register\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08927__B2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 top.DUT.register\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold675 top.DUT.register\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 top.DUT.register\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 top.DUT.register\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _04060_ net456 net535 _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__o211a_2
X_08917_ net279 _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nand2_1
X_09897_ _03937_ net457 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_96_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10004__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _03058_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _03132_ net459 _03868_ net470 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a22o_1
XANTENNA__10939__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ net162 net1535 net413 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11790_ _05620_ _05629_ net130 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__nand3b_1
XANTENNA__07115__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ net175 net1793 net415 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13460_ clknet_leaf_96_clk _01006_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12219__A2_N _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ net188 net1420 net418 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12411_ clknet_leaf_54_clk top.ru.next_FetchedData\[6\] net1077 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10674__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ clknet_leaf_25_clk _00937_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07969__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ top.pad.button_control.debounce top.pad.button_control.noisy vssd1 vssd1
+ vccd1 vccd1 _06131_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ top.lcd.cnt_20ms\[7\] top.lcd.cnt_20ms\[6\] _06074_ vssd1 vssd1 vccd1 vccd1
+ _06090_ sky130_fd_sc_hd__and3_1
XANTENNA__06641__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__A1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ top.a1.data\[11\] net797 _05050_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_56_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ net923 net1395 net875 _05077_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ net177 net2132 net387 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux2_1
XANTENNA__13511__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11086_ net99 net886 net849 net1299 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10489__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10037_ net172 net2261 net530 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
XANTENNA__07354__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10849__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07290__Y _02407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ _05845_ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13727_ clknet_leaf_63_clk _01257_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ net2269 net175 net486 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13658_ clknet_leaf_88_clk _01199_ net1016 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ clknet_leaf_45_clk _00155_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10584__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13589_ clknet_leaf_55_clk _01130_ net1097 vssd1 vssd1 vccd1 vccd1 top.ramload\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_170_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09096__D _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout407 net409 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_8
X_09820_ _04192_ _04816_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__or3_1
Xfanout418 _04994_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
Xfanout429 _04990_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07593__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _03548_ net456 net535 _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__o211a_1
X_06963_ top.DUT.register\[15\]\[21\] net805 net801 top.DUT.register\[31\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_78_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08702_ net1316 net858 net836 _03801_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__a22o_1
X_09682_ _04698_ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__nor2_1
X_06894_ top.DUT.register\[12\]\[24\] net736 net713 top.DUT.register\[25\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XANTENNA__07345__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08633_ _03734_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06699__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10759__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08564_ net902 top.pc\[11\] net537 _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a22o_1
X_07515_ top.DUT.register\[30\]\[14\] net695 net643 top.DUT.register\[10\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
X_08495_ net904 top.pc\[8\] net539 _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a22o_1
XANTENNA__08845__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_A _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06257__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07446_ _02551_ _02559_ _02562_ _02557_ _02550_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__o311a_1
XANTENNA__06320__A1 top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10494__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06871__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ top.DUT.register\[13\]\[4\] net790 net590 top.DUT.register\[20\]\[4\] _02493_
+ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09116_ _04102_ _04113_ _04168_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__or3b_4
X_06328_ _01333_ _01334_ _01335_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__and3b_1
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09047_ _03900_ _03921_ _03940_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__and4b_1
XFILLER_0_130_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06259_ top.ramload\[17\] net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[17\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09022__B1 _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 top.DUT.register\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold461 top.DUT.register\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 top.DUT.register\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold483 top.DUT.register\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 top.DUT.register\[15\]\[17\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_2
Xfanout952 net959 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_2
X_09949_ top.pc\[29\] _04643_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nor2_1
Xfanout963 net969 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_69_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08128__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net978 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09325__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 net994 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_4
X_12960_ clknet_leaf_13_clk _00506_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_129_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 top.DUT.register\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _05737_ _05771_ _05762_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a21o_1
Xhold1161 top.DUT.register\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 top.DUT.register\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07887__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1183 top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10669__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ clknet_leaf_5_clk _00437_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1194 top.DUT.register\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_11842_ _05700_ _05701_ _05696_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_169_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09089__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11773_ _05568_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13512_ clknet_leaf_31_clk _01058_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ net251 top.DUT.register\[24\]\[5\] net416 vssd1 vssd1 vccd1 vccd1 _00863_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__A _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13443_ clknet_leaf_32_clk _00989_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09478__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06862__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ net258 net1742 net420 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13374_ clknet_leaf_38_clk _00920_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload17 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__bufinv_16
Xclkload28 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_4
X_10586_ net617 _04966_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload39 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_58_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12325_ top.lcd.cnt_500hz\[10\] _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ _06075_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__nor2_2
XANTENNA__09013__B1 _02637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11207_ net908 net405 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12187_ _06045_ _06046_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_207_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11138_ net43 net880 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__and2_1
XANTENNA__08119__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__Q top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__B _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11069_ net16 net863 net835 net1192 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_0_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11123__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07327__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10579__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_clk_X clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07300_ top.DUT.register\[14\]\[1\] net795 net728 top.DUT.register\[10\]\[1\] _02416_
+ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a221o_1
XANTENNA__10634__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08280_ net287 _03394_ _03393_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_82_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07231_ top.DUT.register\[17\]\[8\] net776 net582 top.DUT.register\[4\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06853__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07189__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__X _04941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07162_ top.DUT.register\[28\]\[12\] net738 net592 top.DUT.register\[8\]\[12\] _02268_
+ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ top.DUT.register\[13\]\[15\] net790 net774 top.DUT.register\[2\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13433__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__C _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 _04814_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_1
Xfanout215 _04795_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07566__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ _04798_ _04801_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__xnor2_1
Xfanout237 _04762_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
XANTENNA__07030__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _05400_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
X_07995_ top.DUT.register\[25\]\[21\] net637 net633 top.DUT.register\[27\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a22o_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout385_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ top.a1.dataIn\[2\] net813 net457 _04745_ vssd1 vssd1 vccd1 vccd1 _04746_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06946_ top.DUT.register\[13\]\[22\] net789 net723 top.DUT.register\[16\]\[22\] _02062_
+ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07318__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__A _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _04190_ _04679_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__and2b_1
XANTENNA__10489__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ top.DUT.register\[15\]\[25\] net807 net803 top.DUT.register\[31\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout552_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08616_ net278 _03526_ _03530_ net269 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09596_ _01874_ _01877_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08547_ net274 _03429_ _03436_ _02203_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout817_A _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__A _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _02199_ net270 _02370_ net278 vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ top.DUT.register\[19\]\[5\] net674 net670 top.DUT.register\[31\]\[5\] _02545_
+ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10440_ net1624 net193 net510 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
XANTENNA__08046__B2 top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09794__A1 _03715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net2005 net202 net430 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
XANTENNA__10952__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _05960_ _05963_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__nor2_1
X_13090_ clknet_leaf_11_clk _00636_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12041_ _05892_ _05894_ _05883_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__a21oi_1
Xhold280 top.DUT.register\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 top.DUT.register\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07557__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net761 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout771 net773 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
Xfanout782 _01537_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_6
XANTENNA__07309__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 _01529_ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
X_12943_ clknet_leaf_20_clk _00489_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10399__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06449__Y _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ clknet_leaf_116_clk _00420_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06178__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11825_ _05683_ _05684_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11756_ _05582_ _05583_ _05612_ _05614_ _05591_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07088__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ net2319 net181 net498 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06835__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11687_ _05503_ _05544_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__xor2_2
XANTENNA__06625__B _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13426_ clknet_leaf_108_clk _00972_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10638_ net191 net2076 net374 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
Xclkload106 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_6
XFILLER_0_153_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08680__X _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12416__Q top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09785__A1 top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap350_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_113_clk _00903_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10862__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ net206 net1485 net503 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07796__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ _01448_ net742 _06110_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_188_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07260__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ clknet_leaf_24_clk _00834_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12239_ net1145 _06055_ net613 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06800_ top.DUT.register\[10\]\[30\] net728 net583 top.DUT.register\[4\]\[30\] _01916_
+ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a221o_1
X_07780_ top.DUT.register\[5\]\[30\] net543 net638 top.DUT.register\[25\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
X_06731_ top.DUT.register\[3\]\[3\] net694 net666 top.DUT.register\[14\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ top.pc\[20\] _04467_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__nor2_1
X_06662_ top.DUT.register\[26\]\[1\] net681 net653 top.DUT.register\[17\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XANTENNA__10102__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ net288 _03353_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09381_ _01415_ _04411_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__nor2_1
X_06593_ _01643_ _01709_ net825 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__mux2_1
XANTENNA__09068__A3 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net315 _03358_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__nor2_1
XANTENNA__07079__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08263_ _03342_ _03378_ net301 vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout133_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ top.DUT.register\[12\]\[9\] net736 net749 top.DUT.register\[1\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_104_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ _03302_ _03309_ net295 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__mux2_1
XANTENNA__08590__X _03695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07145_ top.DUT.register\[6\]\[13\] net596 net580 top.DUT.register\[4\]\[13\] _02261_
+ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a221o_1
XANTENNA__10772__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1042_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07076_ top.DUT.register\[29\]\[16\] net784 net592 top.DUT.register\[8\]\[16\] _02192_
+ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07539__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07003__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07978_ top.DUT.register\[13\]\[18\] net675 net548 top.DUT.register\[4\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09717_ top.a1.instruction\[8\] _04730_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06929_ _02031_ _02033_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net137 _04667_ _04671_ net823 _04663_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__o221a_1
XFILLER_0_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09665__A_N _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _05438_ net207 vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__nand2_1
XANTENNA__08267__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12590_ clknet_leaf_93_clk _00136_ net998 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08267__B2 _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__A1_N net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11541_ _01395_ _05386_ net248 vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06817__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _05299_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07490__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ clknet_leaf_5_clk _00757_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10423_ net1675 net261 net512 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10682__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13142_ clknet_leaf_104_clk _00688_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _04181_ net615 _04731_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3_1
XANTENNA__10254__Y _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13073_ clknet_leaf_8_clk _00619_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ net144 top.DUT.register\[10\]\[30\] net437 vssd1 vssd1 vccd1 vccd1 _00440_
+ sky130_fd_sc_hd__mux2_1
X_12024_ _05879_ _05882_ _05856_ _05869_ _05871_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_131_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07950__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06179__Y _01400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ clknet_leaf_37_clk _00472_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10857__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ clknet_leaf_59_clk _00403_ net1103 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06907__Y _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ _05658_ _05660_ _05667_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_140_Left_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12788_ clknet_leaf_99_clk _00334_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11739_ _05569_ _05580_ _05555_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06808__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07481__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10592__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_46_clk _00955_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07233__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08950_ net461 _04025_ _04037_ net465 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07901_ _03011_ _03013_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_168_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ net475 _02979_ _02981_ net398 _03928_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_4_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07832_ top.DUT.register\[4\]\[28\] net550 net542 top.DUT.register\[5\]\[28\] _02948_
+ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a221o_1
XFILLER_0_209_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09024__A2_N _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ net356 _02878_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09502_ top.pc\[23\] _04529_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06714_ net826 _01808_ _01829_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__o21ai_4
X_07694_ top.DUT.register\[5\]\[12\] net540 net647 top.DUT.register\[12\]\[12\] _02810_
+ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04467_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__or2_1
X_06645_ top.DUT.register\[23\]\[2\] net565 net641 top.DUT.register\[9\]\[2\] _01761_
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout250_A _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ top.pc\[15\] _04391_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__nand2_1
X_06576_ top.DUT.register\[28\]\[0\] net656 net541 top.DUT.register\[5\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08315_ _03427_ _03428_ net295 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09295_ _04337_ _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08246_ _03359_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08177_ net905 top.pc\[0\] _03290_ net538 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07128_ net322 _02243_ _02224_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06281__A top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07224__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ net325 _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nor2_1
XANTENNA__10007__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10070_ net184 net2142 net446 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07932__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ clknet_leaf_65_clk _01285_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ net1409 net176 net482 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XANTENNA__08495__X _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12711_ clknet_leaf_50_clk _00257_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10677__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ clknet_leaf_79_clk _00006_ net1088 vssd1 vssd1 vccd1 vccd1 top.ru.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ clknet_leaf_12_clk _00188_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ clknet_leaf_60_clk _00119_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11524_ top.a1.dataIn\[16\] _05363_ _05364_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__and3_1
XANTENNA__07463__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06671__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ _05314_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ net1464 net191 net513 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08412__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07215__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11386_ _05234_ _05236_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_185_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13125_ clknet_leaf_39_clk _00671_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ net1626 net203 net519 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
X_13056_ clknet_leaf_12_clk _00602_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ net215 net2013 net434 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__mux2_1
X_12007_ _05864_ _05845_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__and2b_2
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ net217 net1970 net438 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XANTENNA__07923__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A1_N net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ clknet_leaf_113_clk _00455_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10587__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06430_ top.DUT.register\[10\]\[0\] net727 net725 top.DUT.register\[16\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06361_ top.a1.instruction\[6\] _01483_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08100_ _03210_ _03212_ _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__or3_1
XFILLER_0_173_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _03493_ _03542_ _03559_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07454__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06292_ net2328 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[18\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Right_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08031_ top.DUT.register\[22\]\[19\] net552 net628 top.DUT.register\[29\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06662__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold802 top.DUT.register\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07206__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 top.DUT.register\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 top.DUT.register\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 top.DUT.register\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 top.DUT.register\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 top.ramaddr\[30\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold868 top.DUT.register\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ net257 net1733 net451 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__mux2_1
Xhold879 top.DUT.register\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ _04020_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _03937_ _03954_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1005_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nand2_2
XANTENNA__11166__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ net475 _03229_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07746_ top.DUT.register\[12\]\[31\] net650 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__and2_1
XFILLER_0_211_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07677_ _02787_ _02789_ _02791_ _02793_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__or4_1
XANTENNA__10497__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09416_ top.pc\[18\] _04435_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__xnor2_1
X_06628_ _01719_ _01744_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07693__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09347_ _04386_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__and2b_1
XFILLER_0_164_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06559_ top.a1.instruction\[20\] top.a1.instruction\[21\] top.a1.instruction\[24\]
+ _01644_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_101_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ _04305_ _04308_ _04307_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06563__X _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08229_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__nand2_1
XANTENNA__06653__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11240_ _05120_ net1312 net402 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
XANTENNA__09874__X _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08945__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net924 net1294 net876 _05085_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a31o_1
X_10122_ net253 net1565 net444 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ net267 net1677 net448 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07905__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ clknet_leaf_72_clk _01337_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06738__X _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13743_ clknet_leaf_68_clk _01268_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfxtp_1
X_10955_ net1342 net249 net483 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10200__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07684__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08881__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ clknet_leaf_89_clk _01215_ net1013 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
X_10886_ net1680 net259 net407 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08881__B2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06892__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ clknet_leaf_7_clk _00171_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ clknet_leaf_85_clk _00102_ net1020 vssd1 vssd1 vccd1 vccd1 top.pc\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06644__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ _05363_ _05364_ _05334_ _05337_ _05351_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07729__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ clknet_leaf_89_clk _00034_ net1012 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold109 top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11438_ _05265_ _05297_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10870__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11369_ _05220_ _05222_ _05226_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_210_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13108_ clknet_leaf_108_clk _00654_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ clknet_leaf_21_clk _00585_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_198_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07600_ _02223_ _02715_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__and2_1
X_08580_ _03401_ _03573_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_105_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09649__B1 _04224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07531_ top.DUT.register\[15\]\[13\] net687 net627 top.DUT.register\[29\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
XANTENNA__09113__A2 _04163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12554__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ top.DUT.register\[5\]\[6\] net542 net654 top.DUT.register\[17\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XANTENNA__10110__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07675__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09201_ net137 _04247_ _04251_ net918 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_33_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06413_ net809 _01518_ _01528_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__and3_1
XANTENNA__06883__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13040__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07393_ _02470_ _02509_ net313 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09009__A1_N _02795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ top.a1.instruction\[24\] top.a1.instruction\[25\] top.a1.instruction\[26\]
+ top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__and4_1
X_06344_ _01459_ _01462_ _01469_ _01475_ _01461_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a32o_1
XANTENNA__07427__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06824__A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ _03493_ _03883_ _03535_ _03786_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__or4b_1
X_06275_ net1759 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[1\] sky130_fd_sc_hd__and2_1
XANTENNA_fanout213_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ _02089_ _03127_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold610 top.DUT.register\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 top.DUT.register\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold632 top.DUT.register\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 top.lcd.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08927__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 top.DUT.register\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10780__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 top.DUT.register\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top.DUT.register\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__A _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 top.DUT.register\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 top.DUT.register\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09965_ _04191_ _04946_ _04947_ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout582_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _03924_ _04004_ net294 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09896_ net170 top.DUT.register\[1\]\[23\] net390 vssd1 vssd1 vccd1 vccd1 _00145_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _03920_ _03032_ _03029_ _02024_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout847_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ net398 _03128_ _03129_ net475 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__o22a_1
XANTENNA__06558__X _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07729_ net281 net342 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08312__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ net182 net1859 net415 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XANTENNA__10020__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07666__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06874__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ net193 net1726 net419 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ clknet_leaf_54_clk top.ru.next_FetchedData\[5\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_95_clk _00936_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ net920 net118 _06129_ net2221 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__a22o_1
XANTENNA__06626__B1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12272_ top.lcd.cnt_20ms\[6\] _06074_ top.lcd.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ _06089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12175__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11223_ net1262 net404 net369 _05112_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10690__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net52 net880 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10105_ net181 net2119 net387 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__mux2_1
X_11085_ net98 net882 net848 net1263 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ net174 net1803 net530 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
XANTENNA__09343__A2 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_X net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ _05846_ _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ clknet_leaf_63_clk _01256_ net1106 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_193_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ net1523 net179 net486 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12419__Q top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10865__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ net1493 net192 net489 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__mux2_1
X_13657_ clknet_leaf_88_clk _01198_ net1017 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ clknet_leaf_13_clk _00154_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13588_ clknet_leaf_55_clk _01129_ net1097 vssd1 vssd1 vccd1 vccd1 top.ramload\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08606__B2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08082__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ clknet_leaf_80_clk _00085_ net1081 vssd1 vssd1 vccd1 vccd1 top.pc\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12433__RESET_B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09567__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09166__S _04169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07042__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_8
Xfanout419 _04994_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
X_06962_ _02072_ _02074_ _02076_ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__or4_2
XANTENNA__10105__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ top.pc\[6\] net817 net457 _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a211o_1
X_08701_ net902 top.pc\[17\] net537 _03800_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a22o_1
X_09681_ top.pad.keyCode\[1\] top.pad.keyCode\[0\] top.pad.keyCode\[3\] top.pad.keyCode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__or4b_2
X_06893_ top.DUT.register\[29\]\[24\] net786 net732 top.DUT.register\[23\]\[24\] _02009_
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a221o_1
XANTENNA__08542__B1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _02642_ _03733_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nand2_1
XANTENNA__07896__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ net463 _03649_ _03652_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07514_ top.DUT.register\[8\]\[14\] net556 net667 top.DUT.register\[31\]\[14\] _02630_
+ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ net462 _03586_ _03602_ net464 _03599_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08845__A1 top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08845__B2 _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07445_ _02560_ _02561_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__nor2_2
XANTENNA__06856__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10775__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__B _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06320__A2 _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ top.DUT.register\[22\]\[4\] net607 net595 top.DUT.register\[8\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ _02515_ _03357_ _04134_ _04147_ _04167_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__o311a_1
X_06327_ _01461_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08073__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09046_ _03841_ _03865_ _03882_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__and4_1
XANTENNA__07937__X _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07281__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06258_ net1348 net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[16\] sky130_fd_sc_hd__and2_1
XFILLER_0_20_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07820__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold440 top.DUT.register\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09022__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06189_ top.pc\[2\] vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XANTENNA__06560__Y _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 top.DUT.register\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 top.DUT.register\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 top.DUT.register\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 top.DUT.register\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A2 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 top.DUT.register\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 _01419_ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_2
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10015__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout942 net960 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_2
X_09948_ _04928_ _04929_ _04926_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a21oi_1
Xfanout953 net959 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
Xfanout964 net969 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_2
Xfanout975 net978 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_2
Xfanout986 net993 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09325__A2 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net998 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__buf_2
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _04859_ _04861_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 top.DUT.register\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 top.DUT.register\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net125 _05759_ _05770_ _05735_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a22o_1
Xhold1162 top.DUT.register\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 top.DUT.register\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07887__A2 _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ clknet_leaf_20_clk _00436_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_187_Left_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1184 top.DUT.register\[30\]\[6\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 top.DUT.register\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09105__A _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11841_ _05700_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13623__Q net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11772_ _05597_ _05604_ _05614_ _05599_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__o31a_1
XANTENNA__07639__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13511_ clknet_leaf_49_clk _01057_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06847__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ net256 net1816 net416 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10654_ net263 net2079 net420 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__mux2_1
X_13442_ clknet_leaf_11_clk _00988_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__C1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13373_ clknet_leaf_119_clk _00919_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10585_ net141 net1592 net503 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__mux2_1
Xclkload18 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload29 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_4
X_12324_ _06120_ net742 _06119_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_58_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12255_ _06076_ _06077_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__or3_1
XANTENNA__09013__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ net909 top.a1.state\[0\] _05095_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__or3_1
XANTENNA__07024__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12186_ _06037_ _06040_ _06041_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11137_ net922 net1421 net874 _05068_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13732__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ net15 net851 net850 top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08838__B _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net251 net2122 net532 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__mux2_1
XANTENNA__07878__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ clknet_leaf_66_clk _01239_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06838__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10595__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07230_ net297 _02346_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ top.DUT.register\[13\]\[12\] net788 net766 top.DUT.register\[11\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a22o_1
XANTENNA__08055__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07189__B _02305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07263__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ top.DUT.register\[29\]\[15\] net786 net721 top.DUT.register\[26\]\[15\] _02208_
+ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a221o_1
XANTENNA__07802__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09004__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _04814_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
XFILLER_0_10_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_2
Xfanout227 _04778_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_1
X_09802_ _04801_ _04798_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and2b_1
Xfanout238 _04762_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
Xfanout249 _04756_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
X_07994_ top.DUT.register\[31\]\[21\] net668 net541 top.DUT.register\[5\]\[21\] _03110_
+ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06945_ top.DUT.register\[23\]\[22\] net731 net767 top.DUT.register\[11\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a22o_1
X_09733_ _04171_ net817 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout378_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__inv_2
X_06876_ _01986_ _01988_ _01990_ _01992_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__or4_4
XANTENNA__07869__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ _02642_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_2_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09595_ net840 _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout545_A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06268__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net464 _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nor2_1
XANTENNA__08818__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06829__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08477_ _03584_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout712_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07428_ top.DUT.register\[29\]\[5\] net630 net626 top.DUT.register\[16\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07359_ top.DUT.register\[18\]\[5\] net779 net721 top.DUT.register\[26\]\[5\] _02475_
+ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08046__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09243__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11050__A1 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09794__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ net1494 net206 net432 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
X_09029_ _02900_ _04083_ net1162 net890 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_130_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _05878_ _05899_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__xor2_4
XANTENNA__07006__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 top.DUT.register\[31\]\[22\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold281 top.DUT.register\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 top.DUT.register\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout750 net751 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_4
Xfanout761 net763 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_195_Left_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout783 _01537_ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_4
Xfanout794 _01529_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12942_ clknet_leaf_92_clk _00488_ net997 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_27_clk _00419_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _05647_ _05679_ _05643_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11755_ _05612_ _05614_ _05591_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09482__B2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10706_ net1394 net185 net498 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11686_ top.a1.dataIn\[10\] _05544_ _05545_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13425_ clknet_leaf_7_clk _00971_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ net197 net2066 net375 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
Xclkload107 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__inv_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07245__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__B2 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10568_ net209 net1453 net501 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__mux2_1
X_13356_ clknet_leaf_2_clk _00902_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09785__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ _01405_ _01446_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_188_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07737__B _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ net220 net2214 net379 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
X_13287_ clknet_leaf_52_clk _00833_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12238_ net1144 _06063_ net613 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
X_12169_ _06013_ _06018_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_207_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire346_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06771__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
X_06730_ top.DUT.register\[7\]\[3\] net574 net657 top.DUT.register\[28\]\[3\] _01846_
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06661_ net854 _01777_ _01776_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_210_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _02841_ _03371_ _03510_ net472 _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o221a_1
X_09380_ _04405_ _04406_ _04404_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__o21ai_2
X_06592_ _01682_ _01708_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__nor2_2
X_08331_ net476 _02846_ _02849_ net458 _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07484__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07213_ top.DUT.register\[6\]\[9\] net598 net590 top.DUT.register\[20\]\[9\] _02329_
+ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a221o_1
X_08193_ _03305_ _03308_ net320 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__mux2_1
XANTENNA__08028__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07144_ top.DUT.register\[30\]\[13\] net760 net752 top.DUT.register\[17\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a22o_1
XANTENNA__07236__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ top.DUT.register\[13\]\[16\] net788 net730 top.DUT.register\[23\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a22o_1
XANTENNA__10791__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A _04999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__Y _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_A _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ top.DUT.register\[6\]\[18\] net576 net671 top.DUT.register\[19\]\[18\] _03093_
+ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a221o_1
XFILLER_0_199_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09716_ top.a1.instruction\[7\] net744 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nand2_1
X_06928_ top.DUT.register\[19\]\[23\] net750 _02029_ _02044_ vssd1 vssd1 vccd1 vccd1
+ _02045_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04668_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06859_ top.DUT.register\[28\]\[26\] net739 net771 top.DUT.register\[27\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ net840 _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__nor2_4
X_08529_ _03414_ _03635_ net281 vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07475__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _01395_ net248 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08019__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11471_ _05302_ _05331_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__nor2_1
XANTENNA__10963__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09216__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10422_ net1450 net240 net509 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
X_13210_ clknet_leaf_19_clk _00756_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07227__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__A _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06742__A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08975__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ clknet_leaf_103_clk _00687_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10353_ net1500 net139 net519 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13072_ clknet_leaf_114_clk _00618_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10284_ net149 net2273 net434 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__mux2_1
X_12023_ _05872_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__nor2_1
XANTENNA__07573__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout580 net581 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_4
XANTENNA__06753__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout591 _01563_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_4
XANTENNA__10203__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_X net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ clknet_leaf_120_clk _00471_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_33_clk _00402_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11807_ _05661_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_157_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ clknet_leaf_108_clk _00333_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _05554_ _05566_ _05579_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10873__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ _05501_ _05504_ _05528_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13408_ clknet_leaf_12_clk _00954_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07218__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__B2 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13339_ clknet_leaf_1_clk _00885_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__B1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ top.DUT.register\[3\]\[24\] net694 _03014_ _03016_ vssd1 vssd1 vccd1 vccd1
+ _03017_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_168_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ net275 _03400_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nor2_1
XANTENNA__08579__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ top.DUT.register\[1\]\[28\] net705 net673 top.DUT.register\[19\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a22o_1
XANTENNA__06744__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ net356 _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09501_ net917 top.pc\[22\] _04533_ net911 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__o211a_1
X_06713_ net826 _01808_ _01829_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__o21a_1
X_07693_ top.DUT.register\[2\]\[12\] net683 net679 top.DUT.register\[26\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09432_ top.pc\[18\] _04435_ top.pc\[19\] vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a21oi_1
X_06644_ top.DUT.register\[8\]\[2\] net558 net657 top.DUT.register\[28\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ top.pc\[15\] _04391_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__nor2_1
X_06575_ _01646_ _01649_ _01653_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__and3_4
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09446__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout243_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _03301_ _03305_ net320 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XANTENNA__07457__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ top.pc\[11\] _02775_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ net292 _01855_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10783__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout410_A _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08176_ _01501_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07127_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07058_ _02174_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout877_A _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06983__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__B _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__Y _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net1550 net181 net482 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XANTENNA__10958__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12710_ clknet_leaf_46_clk _00256_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11643__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ clknet_leaf_79_clk _00011_ net1085 vssd1 vssd1 vccd1 vccd1 top.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06737__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ clknet_leaf_42_clk _00187_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ clknet_leaf_60_clk _00118_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _05363_ _05364_ top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10693__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11454_ _05268_ _05309_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ net1691 net198 net514 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__mux2_1
X_11385_ _05240_ _05244_ _05238_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_185_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13124_ clknet_leaf_31_clk _00670_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10336_ net2050 net208 net517 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
XANTENNA__07620__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13055_ clknet_leaf_32_clk _00601_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10267_ _04788_ net1849 net434 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__mux2_1
X_12006_ _05860_ _05862_ _05866_ _05837_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__o2bb2a_1
X_10198_ net219 net2106 net439 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07687__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ clknet_leaf_3_clk _00454_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07151__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12839_ clknet_leaf_44_clk _00385_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09428__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06360_ top.a1.instruction\[2\] top.a1.instruction\[3\] _01481_ vssd1 vssd1 vccd1
+ vccd1 _01483_ sky130_fd_sc_hd__or3_2
XANTENNA__07439__B1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06291_ top.ramload\[17\] net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[17\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08030_ top.DUT.register\[7\]\[19\] net572 net656 top.DUT.register\[28\]\[19\] _03146_
+ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_79_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold803 top.DUT.register\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold814 top.DUT.register\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10108__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold825 top.DUT.register\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 top.DUT.register\[13\]\[22\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold847 top.DUT.register\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold858 top.DUT.register\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ net261 net1899 net452 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__mux2_1
Xhold869 top.DUT.register\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _03996_ _04019_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__nand2_1
X_08863_ _03937_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__inv_2
X_08794_ _01746_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__nor2_1
XANTENNA__07390__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ top.DUT.register\[23\]\[31\] net566 net661 top.DUT.register\[18\]\[31\] _02861_
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a221o_1
XANTENNA__10778__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout458_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07676_ top.DUT.register\[7\]\[10\] net572 net647 top.DUT.register\[12\]\[10\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07142__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09415_ _04450_ _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__a21oi_1
X_06627_ _01721_ _01727_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_36_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06276__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ top.pc\[14\] _04378_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or2_1
X_06558_ net747 _01647_ _01658_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__and3_4
XANTENNA__08772__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ _04320_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__or2_1
X_06489_ _01490_ _01498_ _01596_ _01597_ _01605_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09807__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08228_ net298 net354 vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout994_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ _02718_ _02851_ _02857_ _02858_ _03259_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a41o_1
XANTENNA__10018__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11170_ net60 net882 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and2_1
XANTENNA__08711__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net267 net1987 net444 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__mux2_1
XANTENNA__06956__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10052_ net257 net2324 net447 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
XANTENNA__08012__A _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06708__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12551__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ clknet_leaf_72_clk _01336_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10688__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ clknet_leaf_67_clk _01267_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07669__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ net1576 net255 net483 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XANTENNA__07133__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13673_ clknet_leaf_90_clk _01214_ net1012 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
X_10885_ top.DUT.register\[29\]\[1\] net262 net408 vssd1 vssd1 vccd1 vccd1 _01019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12624_ clknet_leaf_117_clk _00170_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12555_ clknet_leaf_85_clk _00101_ net1020 vssd1 vssd1 vccd1 vccd1 top.pc\[20\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08094__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09023__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ _05337_ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12486_ clknet_leaf_90_clk _00033_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ _05265_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ top.a1.dataIn\[22\] top.a1.dataIn\[21\] _05224_ top.a1.dataIn\[23\] vssd1
+ vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_210_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06947__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_108_clk _00653_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ net1358 net142 net523 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
X_11299_ top.a1.row2\[41\] _05157_ _05161_ top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1
+ _05169_ sky130_fd_sc_hd__a22o_1
XANTENNA__08149__A1 _01874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ clknet_leaf_97_clk _00584_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10598__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06580__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ top.DUT.register\[14\]\[13\] net663 net655 top.DUT.register\[28\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07124__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07461_ top.DUT.register\[21\]\[6\] net570 net546 top.DUT.register\[24\]\[6\] _02577_
+ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13281__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09200_ _04249_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nand2_1
X_06412_ net809 _01527_ _01528_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__and3_4
XFILLER_0_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07392_ net321 net334 _02490_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06343_ _01471_ _01474_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ net914 net913 _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ net310 _03515_ _03833_ _04034_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a2111o_1
X_06274_ net1210 net899 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[0\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07832__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08013_ _02089_ _03127_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold600 top.DUT.register\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold611 top.DUT.register\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout206_A _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap330 _03078_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_1
Xhold622 top.DUT.register\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 top.DUT.register\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07495__X _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold644 top.DUT.register\[3\]\[31\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 top.DUT.register\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 top.DUT.register\[30\]\[10\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold677 top.DUT.register\[24\]\[4\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 top.DUT.register\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold699 top.DUT.register\[2\]\[31\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _04656_ net360 net328 top.a1.dataIn\[30\] net363 vssd1 vssd1 vccd1 vccd1
+ _04948_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1115_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _03966_ _04003_ net319 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__mux2_1
X_09895_ _03918_ net455 net534 _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout575_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08846_ net1351 net861 net838 _03938_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07363__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ net311 _03509_ _03871_ net274 _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__o221a_1
XANTENNA__06571__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13624__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10301__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _02842_ _02843_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__and2_2
XFILLER_0_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07115__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ _02775_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ net196 net1761 net419 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__mux2_1
XANTENNA__06574__X _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08076__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ top.pc\[13\] _04359_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ _06129_ _06130_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ _01383_ _06075_ _06088_ net1117 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__o211a_1
XANTENNA__10971__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ top.a1.data\[10\] net796 _05047_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ net923 net1322 net874 _05076_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_56_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ net185 net2058 net386 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__mux2_1
X_11084_ net95 net885 net849 net1159 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ net181 net1698 net530 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
XANTENNA__08000__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07354__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10211__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _05781_ _05806_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__xnor2_2
X_13725_ clknet_leaf_63_clk _01255_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ net1517 net183 net485 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ clknet_leaf_75_clk _01197_ net1082 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ net1824 net195 net490 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ clknet_leaf_32_clk _00153_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08067__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13587_ clknet_leaf_55_clk _01128_ net1097 vssd1 vssd1 vccd1 vccd1 top.ramload\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ net210 net1751 net410 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ clknet_leaf_86_clk _00084_ net1019 vssd1 vssd1 vccd1 vccd1 top.pc\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10881__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12469_ clknet_leaf_74_clk top.ru.next_write_i net1088 vssd1 vssd1 vccd1 vccd1 top.Wen
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout409 _05001_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07593__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ top.DUT.register\[21\]\[21\] net610 net765 top.DUT.register\[19\]\[21\] _02077_
+ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ net462 _03785_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o21ai_2
X_09680_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_1
X_06892_ top.DUT.register\[10\]\[24\] net729 net718 top.DUT.register\[9\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XANTENNA__07345__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ _02642_ _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10121__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ net474 _03664_ _03666_ net394 _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07513_ top.DUT.register\[1\]\[14\] net703 net552 top.DUT.register\[22\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
X_08493_ _03600_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout156_A _04923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07444_ net308 net335 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06394__X _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09211__A _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07375_ top.DUT.register\[18\]\[4\] net778 net583 top.DUT.register\[4\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout323_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1065_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06554__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _03286_ _03371_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o21ba_1
X_06326_ net1114 _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07805__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09045_ _03718_ _03803_ _03823_ _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_131_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06257_ net1429 net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[15\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold430 top.DUT.register\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ top.pc\[1\] vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
Xhold441 top.DUT.register\[16\]\[14\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 top.DUT.register\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 top.DUT.register\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold474 top.DUT.register\[26\]\[9\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 top.DUT.register\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 top.DUT.register\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 net911 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07584__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout932 net960 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
X_09947_ net151 net1437 net392 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__mux2_1
Xfanout943 net945 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
Xfanout954 net959 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net969 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 net978 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
Xfanout987 net993 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_2
X_09878_ _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_2
Xhold1130 top.DUT.register\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1141 top.DUT.register\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1152 top.DUT.register\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _01775_ _03851_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand2_1
Xhold1163 top.lcd.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 top.DUT.register\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06544__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 top.DUT.register\[4\]\[2\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 top.DUT.register\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ _05654_ _05697_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10031__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _05597_ _05614_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__or2_1
XANTENNA__10966__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ clknet_leaf_47_clk _01056_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ net267 net2305 net416 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13441_ clknet_leaf_41_clk _00987_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08049__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ net241 net1209 net419 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ clknet_leaf_18_clk _00918_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10584_ net144 net2250 net503 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload19 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_6
X_12323_ top.lcd.cnt_500hz\[9\] _06118_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07576__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ top.lcd.cnt_20ms\[15\] top.lcd.cnt_20ms\[14\] top.lcd.cnt_20ms\[17\] top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__or4bb_1
XANTENNA__09013__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ top.a1.row1\[63\] _05096_ _05106_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_71_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ _06037_ _06040_ _06044_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10206__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11136_ net42 net880 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__and2_1
XANTENNA__11108__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11067_ net14 net863 net835 net1297 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__o22a_1
XANTENNA__09008__A1_N net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__A1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07327__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11123__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ net256 net2246 net531 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13772__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10876__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__B1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _05818_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13708_ clknet_leaf_64_clk _01238_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09031__A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13639_ clknet_leaf_93_clk net1212 net995 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07160_ _02271_ _02273_ _02274_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__or4_1
XFILLER_0_109_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07091_ top.DUT.register\[28\]\[15\] net740 net736 top.DUT.register\[12\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 _04814_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_1
Xfanout217 _04788_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
X_09801_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__or2_1
XANTENNA__07566__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout239 _04762_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_1
X_07993_ top.DUT.register\[20\]\[21\] net561 net648 top.DUT.register\[12\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a22o_1
X_09732_ net264 net1307 net392 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06944_ top.DUT.register\[30\]\[22\] net761 net755 top.DUT.register\[18\]\[22\] _02050_
+ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a221o_1
XANTENNA__07318__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08515__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08515__B2 _03364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _04684_ _04685_ _04674_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a21o_1
X_06875_ top.DUT.register\[23\]\[25\] net732 net591 top.DUT.register\[20\]\[25\] _01991_
+ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout273_A _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _02664_ _03697_ _02665_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_2_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09594_ top.a1.instruction\[28\] net842 net619 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08545_ _02745_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__xor2_1
XANTENNA__10786__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_A _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _02773_ _03583_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07427_ top.DUT.register\[11\]\[5\] net701 net638 top.DUT.register\[25\]\[5\] _02543_
+ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06284__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07358_ top.DUT.register\[10\]\[5\] net728 net763 top.DUT.register\[30\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10389__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06309_ _01405_ _01446_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__or2_1
X_07289_ top.DUT.register\[17\]\[2\] net753 _02391_ _02405_ vssd1 vssd1 vccd1 vccd1
+ _02406_ sky130_fd_sc_hd__a211o_1
X_09028_ _02925_ net620 net1315 net887 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 top.DUT.register\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10026__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 top.DUT.register\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 top.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07557__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 top.DUT.register\[29\]\[28\] vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06765__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_8
Xfanout751 _01581_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
Xfanout762 net763 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout773 _01557_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07309__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout784 _01534_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
Xfanout795 _01529_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_2
X_12941_ clknet_leaf_113_clk _00487_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13634__Q net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ clknet_leaf_26_clk _00418_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07190__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _05680_ _05643_ _05677_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_29_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ _05612_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__and2_1
X_10705_ net1881 net189 net497 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ _05544_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13424_ clknet_leaf_117_clk _00970_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ net200 net1929 net374 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload108 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13355_ clknet_leaf_4_clk _00901_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ net215 net2067 net501 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__mux2_1
X_12306_ _01446_ net742 _06109_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07796__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13286_ clknet_leaf_19_clk _00832_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_188_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10498_ net226 net2263 net378 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ net1177 _06068_ net612 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ _06018_ _06019_ _06013_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06756__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11119_ net925 net1279 net877 _05059_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_207_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ _05897_ _05957_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a21bo_1
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XANTENNA_wire339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06660_ top.a1.instruction\[22\] net824 _01640_ top.a1.instruction\[30\] vssd1 vssd1
+ vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06591_ _01688_ _01694_ _01700_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06656__Y _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ net396 _02847_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08261_ net296 _03376_ _03349_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08681__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13835__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ top.DUT.register\[27\]\[9\] net772 net768 top.DUT.register\[11\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08192_ _03306_ _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07143_ top.DUT.register\[29\]\[13\] net784 net600 top.DUT.register\[5\]\[13\] _02259_
+ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10240__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07074_ top.DUT.register\[16\]\[16\] net723 net580 top.DUT.register\[4\]\[16\] _02178_
+ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a221o_1
XANTENNA__08474__B1_N _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07539__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08736__B2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06747__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ top.DUT.register\[26\]\[18\] net679 net663 top.DUT.register\[14\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09715_ top.a1.instruction\[9\] top.a1.instruction\[10\] net745 vssd1 vssd1 vccd1
+ vccd1 _04729_ sky130_fd_sc_hd__o21a_1
XANTENNA__11185__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06927_ top.DUT.register\[21\]\[23\] net608 net760 top.DUT.register\[30\]\[23\] _02043_
+ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ _01940_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_27_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06858_ top.DUT.register\[7\]\[26\] net708 _01972_ _01974_ vssd1 vssd1 vccd1 vccd1
+ _01975_ sky130_fd_sc_hd__a211o_1
XANTENNA__07172__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09577_ top.a1.instruction\[27\] net841 net618 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a21oi_1
X_06789_ top.DUT.register\[11\]\[30\] net769 net586 top.DUT.register\[24\]\[30\] _01905_
+ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08528_ _03537_ _03634_ net289 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08672__B1 _03772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ net308 net302 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06582__X _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11470_ _05317_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10421_ net617 _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__nor2_4
XANTENNA__07838__B _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07778__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ clknet_leaf_103_clk _00686_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10352_ top.DUT.register\[12\]\[30\] net144 net520 vssd1 vssd1 vccd1 vccd1 _00504_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06986__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13856__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ clknet_leaf_24_clk _00617_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10283_ net152 net2235 net436 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12022_ _05879_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09117__Y _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout570 _01666_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07950__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout581 _01566_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_4
Xfanout592 _01551_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_45_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07860__Y _02977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ clknet_leaf_18_clk _00470_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06757__X _01874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ clknet_leaf_109_clk _00401_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11806_ _05650_ _05662_ _05664_ _05665_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ clknet_leaf_106_clk _00332_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08258__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11737_ _05555_ _05567_ _05580_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12217__A2_N _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _05501_ _05504_ _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13407_ clknet_leaf_23_clk _00953_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ net616 _04968_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__nand2_4
X_11599_ _05422_ _05452_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ clknet_leaf_15_clk _00884_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06977__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13269_ clknet_leaf_100_clk _00815_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08718__A1 _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11286__A top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ top.DUT.register\[6\]\[28\] net578 net558 top.DUT.register\[8\]\[28\] _02946_
+ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07761_ net827 _02877_ _02617_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a21oi_2
X_09500_ net136 _04523_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12051__D_N top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06712_ net828 _01828_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07692_ _02802_ _02804_ _02806_ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__or4_1
XANTENNA__07154__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ top.pc\[18\] top.pc\[19\] _04435_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06643_ top.DUT.register\[6\]\[2\] net577 _01759_ vssd1 vssd1 vccd1 vccd1 _01760_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06901__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ net917 top.pc\[14\] _04402_ net910 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_121_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06319__S _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06574_ _01672_ net799 _01662_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__and3b_1
XFILLER_0_164_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ _03298_ _03339_ net284 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09293_ top.pc\[11\] _02775_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10461__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__X _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net286 _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__or2_1
XANTENNA__07939__A _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ top.d_ready _01487_ _01491_ _01493_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__or4_1
XFILLER_0_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07126_ _02233_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06968__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07057_ _02166_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__nor2_4
XFILLER_0_100_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10304__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ top.DUT.register\[23\]\[20\] net564 net684 top.DUT.register\[2\]\[20\] _03075_
+ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ net2136 net184 net482 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XANTENNA__07145__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ _04652_ _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12757__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ clknet_leaf_12_clk _00186_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ clknet_leaf_60_clk _00117_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10974__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08952__B _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _05341_ _05365_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06671__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _05275_ _05300_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_190_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ net1530 net202 net513 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__mux2_1
X_11384_ _05240_ _05244_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__nand2_1
XANTENNA__06959__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13123_ clknet_leaf_34_clk _00669_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_185_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ net1969 net213 net517 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13054_ clknet_leaf_32_clk _00600_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ net219 top.DUT.register\[10\]\[11\] net434 vssd1 vssd1 vccd1 vccd1 _00421_
+ sky130_fd_sc_hd__mux2_1
X_12005_ _05841_ _05865_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__and2_1
XANTENNA__10214__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10197_ net224 top.DUT.register\[8\]\[10\] net438 vssd1 vssd1 vccd1 vccd1 _00356_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07923__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07136__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ clknet_leaf_4_clk _00453_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12838_ clknet_leaf_48_clk _00384_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_196_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07439__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12769_ clknet_leaf_40_clk _00315_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08636__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06290_ net2348 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[16\] sky130_fd_sc_hd__and2_1
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06662__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold804 top.DUT.register\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 top.DUT.register\[20\]\[0\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 top.lcd.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 top.DUT.register\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold848 top.DUT.register\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ net240 net1950 net451 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__mux2_1
Xhold859 top.DUT.register\[29\]\[10\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ _03996_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08862_ net461 _03940_ _03953_ net466 _03951_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o221a_2
XANTENNA__10124__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ net357 _02926_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08793_ _03538_ _03570_ _03725_ net271 _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout186_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ top.DUT.register\[10\]\[31\] net646 net642 top.DUT.register\[9\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08529__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07675_ top.DUT.register\[15\]\[10\] net687 net623 top.DUT.register\[16\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1095_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ net915 top.pc\[17\] net910 vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__o21ai_1
X_06626_ _01713_ _01733_ _01736_ _01737_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09345_ top.pc\[14\] _04378_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout520_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06557_ top.DUT.register\[23\]\[0\] net564 net561 top.DUT.register\[20\]\[0\] _01671_
+ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a221o_1
XANTENNA__09868__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09276_ top.pc\[9\] _04297_ top.pc\[10\] vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06488_ _01488_ _01604_ _01600_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_43_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ net324 _01878_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__or2_1
XANTENNA__06653__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06292__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _03182_ _03228_ _02068_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__or3b_1
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout987_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ top.DUT.register\[22\]\[14\] net604 net601 top.DUT.register\[5\]\[14\] _02225_
+ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08089_ _02174_ _03203_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__or2_1
X_10120_ net258 net1308 net443 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10051_ net261 net1694 net449 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
XANTENNA__10034__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07366__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07905__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10969__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_69_clk _01335_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07118__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13741_ clknet_leaf_68_clk _01266_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_119_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10953_ net1942 net266 net483 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XANTENNA__08866__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13672_ clknet_leaf_90_clk _01213_ net1012 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
X_10884_ net2148 net242 net407 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12623_ clknet_leaf_23_clk _00169_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06892__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09602__B1_N net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ clknet_leaf_89_clk _00100_ net1014 vssd1 vssd1 vccd1 vccd1 top.pc\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _05363_ _05364_ _05351_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06644__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12485_ clknet_leaf_90_clk _00032_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10209__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11436_ _05293_ _05295_ _05278_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_128_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11367_ _05224_ _05226_ _05227_ _05223_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__o31a_2
XFILLER_0_21_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ clknet_leaf_106_clk _00652_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ net1697 net144 net524 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11298_ top.a1.row1\[17\] _05155_ _05158_ top.a1.row1\[9\] _05167_ vssd1 vssd1 vccd1
+ vccd1 _05168_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_165_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08149__A2 _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13037_ clknet_leaf_114_clk _00583_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ net150 net1857 net383 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__mux2_1
XANTENNA__07357__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07109__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09649__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ top.DUT.register\[19\]\[6\] net673 net649 top.DUT.register\[12\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06411_ top.a1.instruction\[17\] top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1
+ _01528_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06883__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07391_ _02501_ _02504_ _02506_ _02507_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__nor4_1
XFILLER_0_158_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ top.a1.instruction\[7\] top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 _04183_
+ sky130_fd_sc_hd__and2_2
X_06342_ _01333_ _01470_ _01473_ _01459_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10186__Y _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _03721_ _03744_ _03762_ _03815_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__or4b_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10119__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06273_ net1238 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[31\] sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08012_ _02090_ _03127_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06680__X _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 top.DUT.register\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 top.DUT.register\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 top.pad.keyCode\[0\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold634 top.DUT.register\[19\]\[4\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap353 net354 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
Xhold645 top.DUT.register\[16\]\[15\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 top.DUT.register\[31\]\[7\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 top.DUT.register\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07060__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold678 top.DUT.register\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ _04170_ _04651_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__nor2_1
Xhold689 top.DUT.register\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08113__A _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08914_ _01879_ _01962_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__nand2_1
X_09894_ _04880_ _04884_ _04879_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__or3b_1
XANTENNA__07348__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08845_ top.ru.state\[5\] top.pc\[24\] net539 _03937_ vssd1 vssd1 vccd1 vccd1 _03938_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10789__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08776_ net269 _03704_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07727_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06287__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ net856 _02589_ _02774_ _01615_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_45_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06609_ _01722_ _01724_ _01725_ _01599_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06874__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout902_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ top.DUT.register\[7\]\[15\] net574 net669 top.DUT.register\[31\]\[15\] _02705_
+ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07399__A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ _04368_ _04369_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09273__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06626__A2 _01733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _04293_ _04295_ _04294_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10029__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12270_ _01383_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ net1252 net404 net369 _05111_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11152_ net50 net880 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and2_1
XANTENNA__07051__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ net189 net2161 net386 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11083_ net84 net884 net849 net1288 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__a22o_1
XANTENNA__07339__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__A _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10034_ net185 net1941 net529 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__10699__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__X _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ _05815_ _05842_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13724_ clknet_leaf_66_clk _01254_ net1116 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ net1410 net187 net485 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
XANTENNA__07511__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12473__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_193_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10867_ net2113 net199 net489 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13655_ clknet_leaf_75_clk _01196_ net1091 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10287__X _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ clknet_leaf_37_clk _00152_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13586_ clknet_leaf_54_clk _01127_ net1096 vssd1 vssd1 vccd1 vccd1 top.ramload\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ net212 top.DUT.register\[26\]\[13\] net410 vssd1 vssd1 vccd1 vccd1 _00935_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12537_ clknet_leaf_77_clk _00083_ net1081 vssd1 vssd1 vccd1 vccd1 top.pc\[2\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11071__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ clknet_leaf_79_clk top.ru.next_FetchedInstr\[31\] net1085 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[31\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ _05248_ _05255_ _05256_ net478 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__and4_1
X_12399_ clknet_leaf_61_clk net1140 net1107 vssd1 vssd1 vccd1 vccd1 top.edg2.flip2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07042__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06960_ top.DUT.register\[23\]\[21\] net731 net717 top.DUT.register\[9\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_3_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06891_ top.DUT.register\[22\]\[24\] net607 net780 top.DUT.register\[1\]\[24\] _02007_
+ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a221o_1
X_08630_ _03691_ _03732_ _02663_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10402__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ _02745_ net458 _03656_ net469 _03657_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a221o_1
X_07512_ top.DUT.register\[15\]\[14\] net687 net540 top.DUT.register\[5\]\[14\] _02628_
+ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a221o_1
X_08492_ _02773_ _02830_ _03577_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__or3_1
XFILLER_0_187_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07502__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07443_ net308 net335 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06856__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout149_A _04941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ top.DUT.register\[15\]\[4\] net806 net802 top.DUT.register\[31\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _04162_ _04163_ _04164_ _04165_ _04158_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a41o_1
X_06325_ top.lcd.nextState\[5\] top.lcd.currentState\[5\] _01453_ vssd1 vssd1 vccd1
+ vccd1 _01460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ _03761_ _04096_ _03785_ _03741_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07281__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06256_ top.ramload\[14\] net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold420 top.DUT.register\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ top.Wen vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
Xhold431 top.DUT.register\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold442 top.DUT.register\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold453 top.DUT.register\[19\]\[31\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 top.DUT.register\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 top.DUT.register\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout685_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout911 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_4
Xhold497 top.DUT.register\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net924 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_2
X_09946_ _04019_ net455 net534 _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__o211a_2
XFILLER_0_110_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11117__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net958 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net969 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_2
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_2
Xhold1120 top.DUT.register\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ top.pc\[22\] _04525_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout852_A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net993 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 top.DUT.register\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1003 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09730__A1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1142 top.DUT.register\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 top.DUT.register\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _03032_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__xnor2_1
Xhold1164 top.pad.keyCode\[4\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06298__A top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 top.DUT.register\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 top.DUT.register\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ _03105_ _03153_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ _05629_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__nand2_1
XANTENNA__08297__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ net259 net2252 net414 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06847__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ clknet_leaf_13_clk _00986_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ net617 _04970_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__nand2_4
XFILLER_0_193_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09797__A1 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13859__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ clknet_leaf_0_clk _00917_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10583_ net149 net2002 net501 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ top.lcd.cnt_500hz\[9\] _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06761__A _01874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12253_ top.lcd.cnt_20ms\[13\] top.lcd.cnt_20ms\[12\] top.lcd.cnt_20ms\[11\] top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11204_ _01421_ _05105_ _05096_ net868 vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__o211a_1
XANTENNA__07024__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ _06037_ _06040_ _06041_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_71_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ net922 net1359 net874 _05067_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_196_Right_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07980__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11066_ net12 net852 _05054_ net2307 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__a22o_1
X_10017_ net268 net1678 net531 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10222__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ top.a1.dataIn\[5\] net125 net126 vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__and3_1
XANTENNA__09312__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ clknet_leaf_63_clk _01237_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06838__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ net1542 net259 net487 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
X_11899_ net126 vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13638_ clknet_leaf_90_clk _01179_ net1003 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10892__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13569_ clknet_leaf_61_clk top.a1.nextHex\[0\] net1110 vssd1 vssd1 vccd1 vccd1 _01378_
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ top.DUT.register\[10\]\[15\] net728 net598 top.DUT.register\[6\]\[15\] _02206_
+ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a221o_1
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11289__A top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout207 _05465_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_09800_ top.pc\[14\] _04391_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__nor2_1
Xfanout218 _04788_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
X_07992_ top.DUT.register\[4\]\[21\] net550 net641 top.DUT.register\[9\]\[21\] _03108_
+ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a221o_1
Xfanout229 _04775_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08598__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06943_ top.DUT.register\[22\]\[22\] net605 net597 top.DUT.register\[6\]\[22\] _02059_
+ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a221o_1
X_09731_ _03382_ _04737_ net536 _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09745__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ net908 net909 top.a1.state\[0\] _04676_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__or4_1
XANTENNA__10132__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06874_ top.DUT.register\[28\]\[25\] net740 net777 top.DUT.register\[17\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ net1318 net858 net836 _03716_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a22o_1
X_09593_ _04618_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout266_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ _02798_ _03640_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09222__A _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _02773_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__or2_1
XANTENNA__06829__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13482__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ top.DUT.register\[1\]\[5\] net705 net689 top.DUT.register\[15\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09228__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07357_ top.DUT.register\[23\]\[5\] net733 net714 top.DUT.register\[25\]\[5\] _02473_
+ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout600_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__B _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06308_ _01405_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__nor2_1
X_07288_ top.DUT.register\[20\]\[2\] net589 net581 top.DUT.register\[4\]\[2\] _02404_
+ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06462__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09027_ net1341 net889 _02951_ _04082_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06239_ _01441_ _01443_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10307__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07006__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 top.DUT.register\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold261 top.DUT.register\[27\]\[11\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07408__A2_N top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 top.DUT.register\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 top.DUT.register\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top.pad.button_control.r_counter\[11\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 _01526_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07962__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_4
X_09929_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout763 _01565_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout774 net775 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
Xfanout785 _01534_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_2
X_12940_ clknet_leaf_3_clk _00486_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10042__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ clknet_leaf_44_clk _00417_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10977__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _05634_ _05676_ _05640_ net130 vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09132__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _05606_ _05609_ _05613_ _05610_ _05577_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o32a_2
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10704_ net1725 net192 net497 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
X_11684_ top.a1.dataIn\[11\] _05518_ _05536_ _05539_ vssd1 vssd1 vccd1 vccd1 _05545_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_153_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13423_ clknet_leaf_24_clk _00969_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10635_ net205 net2229 net376 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12511__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload109 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__inv_12
XFILLER_0_125_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13354_ clknet_leaf_118_clk _00900_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ _04788_ net1897 net501 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07245__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a21o_1
X_13285_ clknet_leaf_40_clk _00831_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10217__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10497_ net229 net1868 net381 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12236_ net1176 _06066_ net612 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
XANTENNA__11837__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__A2 _03473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _06017_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_9_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07953__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ net62 net885 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and2_1
X_12098_ _05929_ _05956_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_207_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net24 net851 net850 net1947 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a22o_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09170__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10887__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06590_ top.DUT.register\[25\]\[0\] net636 net632 top.DUT.register\[27\]\[0\] _01706_
+ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08130__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _03350_ _03375_ net284 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07484__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08681__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08681__B2 _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07211_ top.DUT.register\[21\]\[9\] net610 net721 top.DUT.register\[26\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08191_ net322 _02326_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_99_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07142_ top.DUT.register\[16\]\[13\] net723 net748 top.DUT.register\[1\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a22o_1
XANTENNA__07236__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07073_ top.DUT.register\[6\]\[16\] net596 _02177_ _02189_ vssd1 vssd1 vccd1 vccd1
+ _02190_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10127__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09933__A1 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07944__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ top.DUT.register\[27\]\[18\] net631 _03089_ _03091_ vssd1 vssd1 vccd1 vccd1
+ _03092_ sky130_fd_sc_hd__a211o_1
XANTENNA__13735__Q top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06926_ top.DUT.register\[23\]\[23\] net730 net715 top.DUT.register\[9\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
X_09714_ top.a1.instruction\[11\] net745 vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10797__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06857_ top.DUT.register\[29\]\[26\] net786 net782 top.DUT.register\[3\]\[26\] _01973_
+ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a221o_1
X_09645_ _01616_ _01640_ top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _04669_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout550_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13663__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09576_ _01982_ _04590_ _04592_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a21oi_1
X_06788_ top.DUT.register\[18\]\[30\] net778 net774 top.DUT.register\[2\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _03593_ _03633_ net313 vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08121__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08458_ net474 net277 _03565_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_172_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07475__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__inv_2
XANTENNA__07678__Y _02795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ _03333_ _03348_ net287 vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09007__A1_N _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ _04181_ _04183_ net744 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand3_2
XANTENNA__07227__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12220__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ net1896 net147 net517 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XANTENNA__08975__A2 _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12545__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ clknet_leaf_92_clk _00616_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10282_ net157 net1985 net434 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__mux2_1
X_12021_ top.a1.dataIn\[4\] _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__nor2_1
XANTENNA__06738__A1 _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout560 _01673_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_8
Xfanout571 _01666_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
Xfanout582 _01566_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_8
Xfanout593 _01551_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_100_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ clknet_leaf_0_clk _00469_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_202_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10500__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ clknet_leaf_102_clk _00400_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ _05664_ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12785_ clknet_leaf_9_clk _00331_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11736_ _05594_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__nand2_1
XANTENNA__07466__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09860__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06674__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _05469_ _05499_ _05526_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__a2bb2o_1
X_13406_ clknet_leaf_38_clk _00952_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07218__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10618_ net142 net1590 net425 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XANTENNA__08206__A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _05430_ _05457_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13337_ clknet_leaf_59_clk _00883_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10549_ net151 net1792 net428 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09736__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13268_ clknet_leaf_108_clk _00814_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08718__A2 _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ _05981_ _05094_ net866 net2299 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07764__B _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ clknet_leaf_24_clk _00745_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07926__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11286__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07760_ _02867_ _02876_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__or2_4
X_06711_ _01818_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07691_ top.DUT.register\[8\]\[12\] net556 net655 top.DUT.register\[28\]\[12\] _02807_
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09430_ net916 top.pc\[18\] _04466_ net910 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__o211a_1
X_06642_ top.DUT.register\[30\]\[2\] net696 net677 top.DUT.register\[13\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a22o_1
XANTENNA__10410__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ net135 _04389_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_121_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06573_ net747 _01647_ _01652_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_121_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08103__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ net1279 net861 net838 _03426_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09292_ _04334_ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
XANTENNA__07457__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06665__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net315 _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout131_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _01494_ _01501_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ _02237_ _02239_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07056_ _02168_ _02170_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__or3_1
XANTENNA__07090__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10652__Y _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07917__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ top.DUT.register\[21\]\[20\] net568 net671 top.DUT.register\[19\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06909_ _02004_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout932_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ net354 _03003_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ top.pc\[30\] _04643_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__xor2_1
XANTENNA__08893__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _04586_ _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ clknet_leaf_60_clk _00116_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09410__A _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ top.a1.dataIn\[16\] _05305_ _05338_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _05306_ _05307_ _05311_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_152_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ net1412 net205 net515 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ top.a1.dataIn\[19\] _05239_ _05242_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__or3_1
X_10334_ net1860 net217 net517 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__mux2_1
X_13122_ clknet_leaf_10_clk _00668_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07620__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13053_ clknet_leaf_1_clk _00599_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ net226 net1930 net434 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07908__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _05850_ _05857_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_167_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ net228 net1649 net440 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout390 _04734_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_6
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_117_clk _00452_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10230__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08884__B2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06895__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ clknet_leaf_40_clk _00383_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08636__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08636__B2 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ clknet_leaf_14_clk _00314_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06647__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _05571_ _05576_ _05578_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a21o_1
X_12699_ clknet_leaf_2_clk _00245_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
XFILLER_0_126_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12454__Q top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08939__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold805 top.DUT.register\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 top.DUT.register\[5\]\[17\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 top.DUT.register\[30\]\[29\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold838 top.d_ready vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 top.DUT.register\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _01729_ _02954_ _04002_ _04018_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__a211o_1
XANTENNA__10405__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ _03058_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__xnor2_1
X_07812_ net357 _02926_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__nand2_1
X_08792_ net272 _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07743_ top.DUT.register\[2\]\[31\] net685 net543 top.DUT.register\[5\]\[31\] _02859_
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout179_A _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ top.DUT.register\[23\]\[10\] net564 net671 top.DUT.register\[19\]\[10\] _02790_
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__a221o_1
XANTENNA__10140__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06625_ _01733_ _01736_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__or2_2
X_09413_ net131 _04437_ net915 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _04373_ _04374_ _04372_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__o21ai_2
X_06556_ _01650_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__nor2_4
XFILLER_0_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_205_Left_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06638__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ top.pc\[9\] top.pc\[10\] _04297_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__and3_1
X_06487_ _01601_ _01603_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout513_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08226_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _03130_ _03271_ _03273_ _03258_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_134_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07108_ top.DUT.register\[23\]\[14\] net731 net588 top.DUT.register\[20\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07063__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _02175_ _03203_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06810__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ top.DUT.register\[9\]\[17\] net716 net757 top.DUT.register\[3\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a22o_1
XANTENNA__10315__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ net242 net2310 net447 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__C _02903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13740_ clknet_leaf_68_clk _01265_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10050__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ net1605 net260 net482 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
XANTENNA__08866__A1 top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06877__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ clknet_leaf_90_clk _01212_ net1011 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
X_10883_ _04181_ net616 _04731_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ clknet_leaf_92_clk _00168_ net997 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09815__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ clknet_leaf_89_clk _00099_ net1014 vssd1 vssd1 vccd1 vccd1 top.pc\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08094__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ _05363_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ clknet_leaf_90_clk _00031_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ net327 _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09139__X _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ top.a1.dataIn\[23\] top.a1.dataIn\[21\] top.a1.dataIn\[20\] top.a1.dataIn\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or4bb_1
XANTENNA__13766__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10317_ net1563 net148 net521 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ clknet_leaf_7_clk _00651_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10225__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ top.a1.row1\[1\] _05154_ _05160_ top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1
+ _05167_ sky130_fd_sc_hd__a22o_1
XANTENNA__08203__B _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__A3 _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ net155 net2184 net382 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__mux2_1
X_13036_ clknet_leaf_3_clk _00582_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10179_ net1353 net151 net528 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_198_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08306__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07106__Y _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08857__B2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_clk_X clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10895__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ net1129 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_201_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06410_ top.a1.instruction\[15\] top.a1.instruction\[16\] net830 vssd1 vssd1 vccd1
+ vccd1 _01527_ sky130_fd_sc_hd__and3b_2
XANTENNA__11580__A top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ top.DUT.register\[6\]\[4\] net598 net759 top.DUT.register\[2\]\[4\] _02492_
+ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06341_ _01333_ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _03602_ _04068_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__and3_1
XANTENNA__07293__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06272_ net1524 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[30\] sky130_fd_sc_hd__and2_1
XANTENNA__07832__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ _02090_ _03127_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold602 top.DUT.register\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 top.DUT.register\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07045__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 top.DUT.register\[6\]\[22\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold635 top.DUT.register\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold646 top.DUT.register\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 top.DUT.register\[13\]\[13\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 top.DUT.register\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 top.DUT.register\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10135__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09962_ _04944_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__xor2_1
X_08913_ net461 _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__nor2_1
X_09893_ _04882_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_209_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A _01774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net399 _03031_ _03936_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21a_2
XANTENNA__07899__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ _03789_ _03870_ net295 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__mux2_1
XANTENNA__06571__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07726_ net292 net339 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06859__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout630_A _01703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ _01777_ _01635_ net400 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06608_ _01388_ _01488_ _01600_ _01716_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__nand4_1
XFILLER_0_165_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07588_ top.DUT.register\[14\]\[15\] net665 net542 top.DUT.register\[5\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ top.pc\[12\] _04334_ top.pc\[13\] vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a21oi_1
X_06539_ top.a1.instruction\[20\] top.a1.instruction\[21\] net799 vssd1 vssd1 vccd1
+ vccd1 _01656_ sky130_fd_sc_hd__and3_2
XFILLER_0_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09273__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08076__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07284__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09258_ _01413_ net853 net873 _04304_ vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_145_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07823__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ net290 _03324_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09189_ top.pc\[2\] top.pc\[3\] top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09025__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11220_ top.a1.data\[9\] net796 _05043_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__o21a_1
XANTENNA__09576__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09597__A_N _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net922 net1331 net875 _05075_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a31o_1
XANTENNA__10045__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net194 net1932 net387 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__mux2_1
X_11082_ net73 net879 net847 net1157 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10033_ net189 net2025 net529 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
XANTENNA__08000__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _05831_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13723_ clknet_leaf_63_clk _01253_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10935_ net1527 net194 net486 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13654_ clknet_leaf_75_clk _01195_ net1083 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
X_10866_ net1620 net203 net491 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12605_ clknet_leaf_120_clk _00151_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08067__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ clknet_leaf_65_clk _01126_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ net218 net2210 net411 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07275__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12536_ clknet_leaf_93_clk _00082_ net947 vssd1 vssd1 vccd1 vccd1 top.ramstore\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11071__B2 top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12467_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[30\] net1087 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[30\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07027__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _05248_ net478 vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__nand2_1
X_12398_ clknet_leaf_60_clk top.edg2.button_i net1100 vssd1 vssd1 vccd1 vccd1 top.edg2.flip1
+ sky130_fd_sc_hd__dfrtp_1
X_11349_ top.a1.row1\[63\] _05140_ _05183_ top.a1.row1\[111\] _05212_ vssd1 vssd1
+ vccd1 vccd1 _05213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09744__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11575__A top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13019_ clknet_leaf_0_clk _00565_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ top.DUT.register\[3\]\[24\] net782 net709 top.DUT.register\[7\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
XANTENNA__09316__Y _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _03653_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__and2_1
X_07511_ top.DUT.register\[7\]\[14\] net572 net675 top.DUT.register\[13\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
X_08491_ _02830_ _03577_ _02773_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_202_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07442_ _02555_ _02556_ _02558_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ net297 _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06324_ top.lcd.nextState\[4\] net845 net843 top.lcd.currentState\[4\] net1114 vssd1
+ vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__o221a_2
XFILLER_0_174_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11062__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _03545_ _03638_ _03689_ _03732_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__and4_1
XANTENNA__07266__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09043_ _03649_ _03672_ _03698_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__or4_1
X_06255_ net1180 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07018__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 top.DUT.register\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06186_ top.Ren vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
Xhold421 top.DUT.register\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold432 top.DUT.register\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08766__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 top.DUT.register\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 top.DUT.register\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 top.DUT.register\[30\]\[17\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13270__RESET_B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 top.DUT.register\[4\]\[11\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 top.DUT.register\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07963__A _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold498 top.DUT.register\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__B2 _01400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _04192_ _04930_ _04925_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__o21ai_1
Xfanout912 top.a1.instruction\[12\] vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout580_A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_147_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout934 net937 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net950 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_2
Xfanout956 net958 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
Xfanout967 net969 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
X_09876_ top.pc\[22\] _04525_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__nand2_1
Xhold1110 top.DUT.register\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout978 net994 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_2
Xhold1121 top.DUT.register\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout989 net993 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1132 top.DUT.register\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _03181_ _03899_ _03182_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a21oi_1
Xhold1143 top.DUT.register\[9\]\[31\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 top.DUT.register\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1165 top.DUT.register\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06544__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1176 top.DUT.register\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 top.DUT.register\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net394 _03842_ _03854_ net474 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a22o_1
Xhold1198 top.DUT.register\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07709_ _02666_ _02695_ _02799_ _02823_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or4_1
X_08689_ _03749_ _03788_ net320 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ net262 top.DUT.register\[24\]\[1\] net416 vssd1 vssd1 vccd1 vccd1 _00859_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_156_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07711__A_N _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08049__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ net141 net1662 net377 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07257__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13370_ clknet_leaf_14_clk _00916_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ net151 net1875 net503 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12321_ _06118_ net742 _06117_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__and3b_1
XFILLER_0_91_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06761__B _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07009__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ top.lcd.cnt_20ms\[9\] top.lcd.cnt_20ms\[7\] top.lcd.cnt_20ms\[6\] top.lcd.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_170_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11203_ _01385_ _01425_ _01427_ _01402_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__o22a_1
X_12183_ _06025_ _06033_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net41 net881 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11065_ net11 net851 net850 net2350 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__a22o_1
XANTENNA__10503__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net257 net1558 net530 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
XANTENNA_input27_X net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _05796_ _05798_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_174_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13706_ clknet_leaf_63_clk _01236_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ net1709 net264 net488 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
X_11898_ _05717_ _05722_ _05748_ _05720_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a22o_1
X_13637_ clknet_leaf_111_clk net1179 net947 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09237__A1 _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10849_ net1833 net139 net496 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ clknet_leaf_62_clk _01114_ net1109 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06952__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09159__A2_N _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07400__X _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08996__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ clknet_leaf_91_clk _00065_ net1003 vssd1 vssd1 vccd1 vccd1 top.ramstore\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13499_ clknet_leaf_0_clk _01045_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_183_Left_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout208 net211 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_2
Xfanout219 _04781_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
X_07991_ top.DUT.register\[11\]\[21\] net701 net546 top.DUT.register\[24\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09730_ top.a1.dataIn\[1\] _01499_ _04740_ top.pc\[1\] _04736_ vssd1 vssd1 vccd1
+ vccd1 _04743_ sky130_fd_sc_hd__a221o_1
XANTENNA__10413__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06942_ top.DUT.register\[28\]\[22\] net739 net748 top.DUT.register\[1\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a22o_1
XANTENNA__06399__A top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__inv_2
X_06873_ top.DUT.register\[12\]\[25\] net736 net714 top.DUT.register\[25\]\[25\] _01989_
+ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ net902 top.pc\[13\] net537 _03715_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__a22o_1
X_09592_ top.pc\[28\] _04606_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__xor2_1
XANTENNA__09503__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ _02745_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout161_A _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout259_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__B _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _02828_ _03550_ _02612_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07425_ top.DUT.register\[21\]\[5\] net570 net634 top.DUT.register\[27\]\[5\] _02541_
+ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1070_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12232__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ top.DUT.register\[28\]\[5\] net740 net780 top.DUT.register\[1\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06307_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__nand3_1
X_07287_ top.DUT.register\[27\]\[2\] net771 net755 top.DUT.register\[18\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06238_ _01443_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__inv_2
X_09026_ net1229 net887 _03002_ net622 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout795_A _01529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06169_ top.edg2.flip2 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
Xhold240 top.DUT.register\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 top.a1.data\[4\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 top.DUT.register\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 top.DUT.register\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 top.DUT.register\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 top.DUT.register\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout962_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _01548_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_4
Xfanout731 net733 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_8
Xfanout742 _06107_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10323__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ top.pc\[27\] _04606_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__and2_1
Xfanout753 _01578_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_4
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08301__B net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 _01556_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
XFILLER_0_204_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout786 _01534_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
Xfanout797 _05010_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _04843_ _04846_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12870_ clknet_leaf_22_clk _00416_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07190__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _05669_ _05673_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_1_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07478__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _05554_ _05570_ _05579_ _05600_ _05562_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_159_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10703_ net1438 net196 net498 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XANTENNA__12547__Q top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ _05518_ _05536_ _05539_ top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 _05544_
+ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_81_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13422_ clknet_leaf_93_clk _00968_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11026__B2 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ net211 net2255 net374 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__B1 _01920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13353_ clknet_leaf_27_clk _00899_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ net221 net1919 net501 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__mux2_1
XANTENNA__06491__B _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ _01445_ net742 _06108_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13284_ clknet_leaf_28_clk _00830_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10496_ net234 net1596 net381 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12235_ net1146 _06065_ net613 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
X_12166_ _05997_ _06007_ _06009_ _06021_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_9_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06756__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ net925 net1340 net877 _05058_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a31o_1
XANTENNA__10233__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _05897_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_207_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08211__B _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ net13 net851 net850 net1759 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a22o_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_204_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12999_ clknet_leaf_56_clk _00545_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12457__Q top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07210_ net321 _02325_ _02306_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12214__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ net322 _02346_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ top.DUT.register\[24\]\[13\] net585 _02246_ _02257_ vssd1 vssd1 vccd1 vccd1
+ _02258_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_191_Left_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10408__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09630__A1 top.a1.instruction\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ top.DUT.register\[5\]\[16\] net600 net588 top.DUT.register\[20\]\[16\] _02188_
+ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a221o_1
XANTENNA__09021__A2_N net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07641__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06747__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10143__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ top.DUT.register\[23\]\[18\] net564 net635 top.DUT.register\[25\]\[18\] _03090_
+ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a221o_1
X_09713_ top.a1.instruction\[11\] net745 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__and2_1
X_06925_ _02035_ _02037_ _02039_ _02041_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_126_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout376_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__A top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _01920_ _04656_ _04658_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06856_ top.DUT.register\[18\]\[26\] net779 net768 top.DUT.register\[11\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07172__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ net136 _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06787_ top.DUT.register\[13\]\[30\] net790 net736 top.DUT.register\[12\]\[30\] _01903_
+ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout543_A _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ net321 _02325_ _02347_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08457_ net476 _02830_ _02833_ net458 _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a221o_1
XFILLER_0_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08672__A2 _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ _01640_ top.a1.instruction\[26\] _01389_ _01615_ vssd1 vssd1 vccd1 vccd1
+ _02525_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12205__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08388_ net269 _03498_ _03499_ net280 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07339_ top.DUT.register\[13\]\[6\] net790 net582 top.DUT.register\[4\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XANTENNA__10318__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10350_ net2149 net150 net518 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XANTENNA__07632__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06986__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _02795_ net620 net1258 net887 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__a2bb2o_1
X_10281_ net160 net2043 net436 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _05830_ _05864_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09408__A _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 _01687_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_8
Xfanout561 _01673_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_4
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_4
Xfanout583 _01566_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
Xfanout594 _01551_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_8
X_12922_ clknet_leaf_15_clk _00468_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07699__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08360__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12853_ clknet_leaf_82_clk _00399_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11804_ _05622_ _05628_ net129 vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12784_ clknet_leaf_115_clk _00330_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11735_ _05555_ _05579_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08193__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ top.a1.dataIn\[12\] _05437_ _05466_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13302__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13405_ clknet_leaf_119_clk _00951_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net143 net2289 net425 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10228__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ _05430_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and2_1
XANTENNA__08206__B _02469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07885__X _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ clknet_leaf_36_clk _00882_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07623__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10548_ net156 net2306 net427 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06977__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ clknet_leaf_95_clk _00813_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10479_ net166 net2187 net507 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12218_ net1261 net866 net831 _05994_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a22o_1
XANTENNA__09318__A _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ clknet_leaf_97_clk _00744_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08222__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ _06007_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09752__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10898__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _01820_ _01822_ _01824_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__or4_1
X_07690_ top.DUT.register\[1\]\[12\] net703 net675 top.DUT.register\[13\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07154__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08351__B2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06641_ top.DUT.register\[11\]\[2\] net700 net636 top.DUT.register\[25\]\[2\] _01757_
+ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a221o_1
XANTENNA__06901__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ net821 _04397_ _04400_ net131 net917 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_121_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06572_ _01659_ _01672_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nor2_4
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08311_ net905 top.pc\[2\] net539 _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09291_ top.pc\[11\] _04320_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__nor2_1
XANTENNA__06683__Y _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _01739_ _03314_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13043__RESET_B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09064__C1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10138__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _03278_ _03286_ _03289_ _02524_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07124_ top.DUT.register\[9\]\[14\] net715 net584 top.DUT.register\[24\]\[14\] _02240_
+ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a221o_1
XANTENNA__07614__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06968__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ top.DUT.register\[27\]\[17\] net771 net589 top.DUT.register\[20\]\[17\] _02171_
+ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1033_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout493_A _04999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ top.DUT.register\[14\]\[20\] net664 net632 top.DUT.register\[27\]\[20\] _03073_
+ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ net324 _02023_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__nand2_1
XANTENNA__13627__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10601__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ net354 _03003_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__and2_1
XANTENNA__07145__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09627_ _04633_ _04635_ _04631_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__o21ai_1
X_06839_ top.DUT.register\[18\]\[27\] net754 _01944_ _01955_ vssd1 vssd1 vccd1 vccd1
+ _01956_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout925_A _01400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A2 _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ top.pc\[26\] _04576_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08509_ net283 _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09489_ _04520_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11520_ _05363_ _05364_ _05342_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_175_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09410__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07853__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11451_ _05306_ _05307_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ net1413 net208 net513 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
XANTENNA__09837__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07605__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11382_ _05239_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06959__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ clknet_leaf_43_clk _00667_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ net1618 net221 net518 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13052_ clknet_leaf_17_clk _00598_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ net230 net2153 net436 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__mux2_1
X_12003_ _05861_ _05863_ _05860_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08030__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10195_ net232 net1518 net440 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_4_13__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout391 _04734_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
XFILLER_0_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10511__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08333__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ clknet_leaf_27_clk _00451_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13554__RESET_B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12836_ clknet_leaf_29_clk _00382_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12767_ clknet_leaf_47_clk _00313_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11718_ _05571_ _05576_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07844__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ clknet_leaf_16_clk _00244_ net989 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__dlymetal6s2s_1
X_11649_ _05422_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
XFILLER_0_126_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold806 top.DUT.register\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold817 top.DUT.register\[21\]\[4\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_52_clk _00865_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold828 top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold839 top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08021__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _03030_ _03930_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08572__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _01898_ _02926_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__nor2_1
XANTENNA__11171__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08791_ _03810_ _03885_ net290 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
XANTENNA__06583__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07742_ top.DUT.register\[13\]\[31\] net677 net625 top.DUT.register\[16\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XANTENNA__09006__A1_N _02610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ top.DUT.register\[26\]\[10\] net679 net552 top.DUT.register\[22\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09412_ net135 _04442_ _04449_ net821 vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o22a_1
XFILLER_0_189_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06624_ _01733_ _01736_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11760__B top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ net915 top.pc\[13\] _04384_ net910 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__o211a_1
X_06555_ top.a1.instruction\[20\] top.a1.instruction\[21\] top.a1.instruction\[24\]
+ net799 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__or4bb_4
XANTENNA__08627__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _04317_ _04318_ _04319_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07835__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06486_ _01388_ top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08225_ _03333_ _03340_ net294 vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout506_A _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08156_ _03082_ _03132_ _03272_ _03260_ _03159_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_134_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07107_ net322 _02223_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08087_ _02175_ _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07038_ _02133_ _02154_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07366__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net356 _02522_ _04074_ net399 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__o211a_1
XFILLER_0_199_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10331__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07118__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ net2035 net261 net484 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13670_ clknet_leaf_90_clk _01211_ net1012 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
X_10882_ net1452 net139 net491 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ clknet_leaf_113_clk _00167_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08079__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09815__A1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12552_ clknet_leaf_84_clk _00098_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[17\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__07826__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08037__A _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ _05323_ _05359_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__xor2_4
X_12483_ clknet_leaf_90_clk _00030_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11434_ _05259_ _05262_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_80_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10506__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_100_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11365_ top.a1.dataIn\[31\] top.a1.dataIn\[25\] top.a1.dataIn\[24\] top.a1.dataIn\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__nand4_1
X_13104_ clknet_leaf_116_clk _00650_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10316_ net2056 net152 net523 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11296_ top.a1.row1\[121\] _05129_ _05136_ top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1
+ _05166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13035_ clknet_leaf_5_clk _00581_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08003__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10247_ net160 net1265 net383 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__mux2_1
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_2
XANTENNA__07357__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09155__X _04208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ net1435 net157 net525 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10241__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07109__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08857__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ net1128 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_202_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12819_ clknet_leaf_110_clk _00365_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13799_ clknet_leaf_69_clk _01324_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06340_ _01458_ _01331_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__and2b_1
XANTENNA__09050__B _03364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07817__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06271_ net1196 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[29\] sky130_fd_sc_hd__and2_1
XFILLER_0_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ net827 _03126_ _02617_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a21o_1
XANTENNA__07786__A _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 top.DUT.register\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 top.DUT.register\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10416__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap333 _02660_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_1
Xhold625 top.DUT.register\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold636 top.DUT.register\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 top.DUT.register\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 top.DUT.register\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _04933_ _04934_ _04935_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__o21a_1
Xhold669 top.a1.row2\[2\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08912_ _02957_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ _04868_ _04873_ _04881_ _04192_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a31o_1
XANTENNA__07348__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08843_ _03368_ _03921_ _03932_ net465 _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout191_A _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10151__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _03824_ _03869_ net317 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07725_ net292 net339 vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout456_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07656_ _02770_ _02771_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nor2_2
XANTENNA__06865__A _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06607_ net912 top.a1.instruction\[14\] _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _02697_ _02699_ _02701_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__or4_1
XFILLER_0_165_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ top.pc\[12\] top.pc\[13\] _04334_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06538_ top.DUT.register\[6\]\[0\] net577 net704 top.DUT.register\[1\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ net137 _04296_ _04299_ net133 _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o221a_1
XFILLER_0_161_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06469_ net809 _01518_ _01536_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _03320_ _03323_ net315 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ top.pc\[2\] top.pc\[3\] top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_78_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08139_ _03253_ _03254_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__nor2_1
XANTENNA__09430__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10326__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11150_ net49 net881 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and2_1
XANTENNA__08784__B2 _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10101_ net196 net1955 net387 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__mux2_1
X_11081_ net72 net877 _01441_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__o21a_1
XANTENNA__08536__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09733__A0 _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07339__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net192 net2238 net529 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
XANTENNA__10061__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__C top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _05842_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__or2_1
XANTENNA__08974__B _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ clknet_leaf_62_clk _01252_ net1106 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ net1604 net197 net486 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07511__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13653_ clknet_leaf_75_clk _01194_ net1084 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
X_10865_ net1391 net210 net489 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ clknet_leaf_18_clk _00150_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13584_ clknet_leaf_65_clk _01125_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10796_ net219 top.DUT.register\[26\]\[11\] net411 vssd1 vssd1 vccd1 vccd1 _00933_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ clknet_leaf_76_clk _00081_ net1082 vssd1 vssd1 vccd1 vccd1 top.ramstore\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08472__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06781__Y _01898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12466_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[29\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[29\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ _05268_ _05273_ _05275_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a211oi_4
XANTENNA__10236__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12397_ _01494_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__inv_2
XANTENNA__08214__B _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ top.a1.row2\[15\] _05188_ _05187_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06786__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ top.lcd.nextState\[5\] top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05150_
+ sky130_fd_sc_hd__nand2b_1
X_13018_ clknet_leaf_16_clk _00564_ net987 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09326__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06538__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09760__S _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07510_ _02620_ _02622_ _02624_ _02626_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__or4_1
X_08490_ net472 _03597_ _03598_ _02522_ _03592_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o221a_1
XANTENNA__06685__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07502__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07441_ net302 net342 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13838__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07372_ _02479_ _02488_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__nor2_4
XFILLER_0_146_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09111_ _03775_ _03804_ _03856_ _03893_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06323_ top.lcd.nextState\[3\] net845 net843 top.lcd.currentState\[3\] net1114 vssd1
+ vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__o221a_2
XTAP_TAPCELL_ROW_118_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06691__Y _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10270__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ _03606_ _04094_ _03626_ _03586_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__or4bb_1
X_06254_ net1197 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[12\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold400 top.DUT.register\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10146__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06185_ top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
Xhold411 top.DUT.register\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 top.DUT.register\[14\]\[1\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08766__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold433 top.DUT.register\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 top.DUT.register\[29\]\[27\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 top.DUT.register\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 top.DUT.register\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold477 top.DUT.register\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07963__B _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout902 net904 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_2
X_09944_ _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold488 top.DUT.register\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
Xhold499 top.DUT.register\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 _01400_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_2
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11117__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net950 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_2
X_09875_ net179 net1758 net391 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__mux2_1
Xhold1100 top.ramload\[8\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout573_A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1111 top.DUT.register\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net982 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 top.DUT.register\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net1346 net858 net836 _03919_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__a22o_1
Xhold1133 top.DUT.register\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1144 top.DUT.register\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 top.DUT.register\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 top.DUT.register\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08757_ _03485_ _03570_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__o21ai_1
Xhold1177 top.DUT.register\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 top.DUT.register\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 top.DUT.register\[21\]\[30\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B _03888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07708_ _02641_ _02720_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__or2_1
XANTENNA__06595__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ _03297_ _03337_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07639_ top.DUT.register\[7\]\[8\] net574 net701 top.DUT.register\[11\]\[8\] _02755_
+ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10650_ net144 net2338 net377 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12539__RESET_B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ top.pc\[12\] _04334_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_24_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ net157 net1579 net501 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__mux2_1
XANTENNA__10261__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[8\] _06115_ vssd1 vssd1 vccd1 vccd1
+ _06118_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10056__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ net2015 _05104_ _05096_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08757__A1 _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ _06037_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06768__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net922 net1344 net874 _05066_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a31o_1
XANTENNA__07980__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net10 net851 net850 top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__a22o_1
X_10015_ net263 net2301 net532 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__mux2_1
XANTENNA__07193__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06940__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06410__A_N top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _05811_ _05812_ _05821_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13705_ clknet_leaf_63_clk _01235_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_10917_ net1404 net240 net486 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
X_11897_ _05745_ _05746_ _05756_ _05754_ _05750_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a311o_1
XFILLER_0_67_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ clknet_leaf_92_clk net1172 net997 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
X_10848_ net1292 net145 net496 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13567_ clknet_leaf_23_clk _01113_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ net154 net2054 net370 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__mux2_1
XANTENNA__06952__B _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12518_ clknet_leaf_111_clk _00064_ net947 vssd1 vssd1 vccd1 vccd1 top.ramstore\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ clknet_leaf_15_clk _01044_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12449_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[12\] net1077 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06471__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_07990_ _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06941_ top.DUT.register\[29\]\[22\] net785 net581 top.DUT.register\[4\]\[22\] _02055_
+ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a221o_1
X_09660_ _04678_ _04679_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__or3_1
X_06872_ top.DUT.register\[26\]\[25\] net721 net709 top.DUT.register\[7\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net463 _03698_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_207_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09591_ _04599_ _04601_ _04598_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _02799_ _03625_ _02326_ _02796_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13660__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08473_ net1293 net860 net837 _03582_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout154_A _04923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07424_ top.DUT.register\[13\]\[5\] net678 net551 top.DUT.register\[4\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12632__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07355_ top.DUT.register\[14\]\[5\] net795 net717 top.DUT.register\[9\]\[5\] _02471_
+ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout321_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06306_ net2302 top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07286_ _02396_ _02398_ _02400_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__or4_1
XANTENNA__06998__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _02977_ net621 net1188 net890 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a2bb2o_1
X_06237_ wb.curr_state\[0\] _01442_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__nand2_1
XANTENNA__06462__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13040__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09936__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 top.DUT.register\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold241 top.DUT.register\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout690_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 top.DUT.register\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 top.DUT.register\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 top.DUT.register\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__A1 top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 top.DUT.register\[28\]\[0\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold296 top.DUT.register\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_X net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout710 _01568_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
Xfanout721 _01548_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_8
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_8
X_09927_ top.pc\[26\] _04590_ _04908_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a21oi_1
Xfanout743 _06107_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_1
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 _01575_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_4
Xfanout765 _01561_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 _01555_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_8
Xfanout787 _01534_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_2
X_09858_ top.pc\[20\] _04494_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__xnor2_1
Xfanout798 _05009_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07175__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ net276 _03556_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21ai_1
X_09789_ _04784_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__nor2_1
XANTENNA__06922__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ _05634_ _05680_ _05677_ _05643_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_1_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _05594_ _05596_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__C top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_166_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ net1619 net202 net497 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11682_ _05501_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_81_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13421_ clknet_leaf_113_clk _00967_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ net212 net2341 net374 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13352_ clknet_leaf_31_clk _00898_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ net226 net2048 net501 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06989__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 _06108_
+ sky130_fd_sc_hd__or2_1
X_13283_ clknet_leaf_34_clk _00829_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10495_ net236 net2049 net380 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
X_12234_ net1143 top.a1.dataIn\[0\] net613 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12165_ top.a1.dataIn\[2\] _06007_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__nor3_1
XANTENNA__10514__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07953__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11116_ net51 net885 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and2_1
XFILLER_0_208_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12096_ _05930_ _05942_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_207_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net2 net862 net834 net1210 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__o22a_1
XANTENNA__13683__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08902__B2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06913__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12998_ clknet_leaf_22_clk _00544_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11949_ _05808_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_71_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08130__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ clknet_leaf_73_clk _01160_ net1120 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07140_ top.DUT.register\[28\]\[13\] net738 net604 top.DUT.register\[22\]\[13\] _02256_
+ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ top.DUT.register\[9\]\[16\] net715 net750 top.DUT.register\[19\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10424__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07944__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ top.DUT.register\[20\]\[18\] net560 net655 top.DUT.register\[28\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a22o_1
X_09712_ net824 _01634_ _01599_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or3b_1
X_06924_ top.DUT.register\[8\]\[23\] net592 net588 top.DUT.register\[20\]\[23\] _02040_
+ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a221o_1
XANTENNA__07157__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09643_ _04665_ _04666_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__xnor2_1
X_06855_ top.DUT.register\[15\]\[26\] net806 net802 top.DUT.register\[31\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a22o_1
XANTENNA__06904__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _04599_ _04601_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__xnor2_1
X_06786_ top.DUT.register\[28\]\[30\] net741 net794 top.DUT.register\[14\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
X_08525_ _02517_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08657__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout536_A _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08456_ net396 _02831_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07321__X _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07407_ _01731_ _01743_ _01859_ _02520_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nand4_2
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _03309_ _03324_ net295 vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07338_ top.DUT.register\[21\]\[6\] net610 net769 top.DUT.register\[11\]\[6\] _02454_
+ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07269_ top.DUT.register\[28\]\[3\] net741 _02372_ _02374_ vssd1 vssd1 vccd1 vccd1
+ _02386_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09008_ net331 net620 net1362 net888 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10280_ net163 net2311 net437 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A2 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_8
Xfanout551 _01687_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
Xfanout562 _01673_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_8
Xfanout573 _01657_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_4
Xfanout584 net585 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 _01551_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09424__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_44_clk _00467_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09143__B _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ clknet_leaf_103_clk _00398_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12558__Q top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11803_ _05628_ net129 _05622_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_14_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12783_ clknet_leaf_21_clk _00329_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11734_ _05549_ _05553_ _05580_ _05551_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a31o_1
XANTENNA__07320__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06674__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ _05497_ _05498_ _05470_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10509__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10616_ net147 net2278 net422 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
X_13404_ clknet_leaf_17_clk _00950_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ _05414_ _05426_ _05434_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13335_ clknet_leaf_112_clk _00881_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07623__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10547_ net158 net1701 net426 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13342__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13266_ clknet_leaf_106_clk _00812_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ net172 net1659 net506 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12217_ _06006_ _05094_ net866 net1931 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10244__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13197_ clknet_leaf_115_clk _00743_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09318__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _05998_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12079_ _05932_ _05933_ _05937_ _05938_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a2111o_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06640_ top.DUT.register\[2\]\[2\] net684 net632 top.DUT.register\[27\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_32_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06571_ top.DUT.register\[14\]\[0\] net664 net549 top.DUT.register\[4\]\[0\] _01685_
+ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_121_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ net394 _03407_ _03424_ net469 _03422_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a221o_2
XANTENNA__08103__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ top.pc\[11\] _04320_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ net303 _03356_ _03326_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__a21o_1
XANTENNA__06665__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10419__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08172_ _01719_ _03288_ _03287_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09064__B1 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ top.DUT.register\[3\]\[14\] net782 net776 top.DUT.register\[17\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07054_ top.DUT.register\[28\]\[17\] net739 net800 top.DUT.register\[31\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__07090__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10154__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1026_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A _05002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ top.DUT.register\[22\]\[20\] net553 net636 top.DUT.register\[25\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a22o_1
X_06907_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07887_ net825 _03002_ _02617_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout653_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07035__Y _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06838_ top.DUT.register\[13\]\[27\] net788 net756 top.DUT.register\[3\]\[27\] _01954_
+ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a221o_1
X_09626_ _04649_ _04650_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ _04569_ _04572_ _04570_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ top.DUT.register\[22\]\[29\] net604 net766 top.DUT.register\[11\]\[29\] _01881_
+ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout820_A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ net307 _01941_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ top.pc\[22\] _04511_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__or2_1
XANTENNA__07302__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ net1295 net860 net838 _03549_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10329__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _05272_ _05296_ _05309_ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_190_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ net1911 net212 net513 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__mux2_1
X_11381_ top.a1.dataIn\[20\] _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120_ clknet_leaf_13_clk _00666_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ net2125 net226 net517 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__mux2_1
XANTENNA__08323__A _01856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13051_ clknet_leaf_1_clk _00597_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10064__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ net232 net2114 net436 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07369__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11165__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _05850_ _05857_ _05838_ _05840_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__a211o_2
XANTENNA__07908__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net238 net2019 net440 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11684__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_6
Xfanout381 _04989_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_8
Xfanout392 _04734_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_6
XFILLER_0_205_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08333__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ clknet_leaf_26_clk _00450_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08993__A _04078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06895__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12835_ clknet_leaf_34_clk _00381_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_26_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12766_ clknet_leaf_39_clk _00312_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07402__A _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _05515_ _05573_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__xnor2_2
XANTENNA__06647__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ clknet_leaf_55_clk _00243_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10239__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ _05453_ _05484_ _05452_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a21bo_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11579_ _05432_ _05433_ _05404_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold807 top.DUT.register\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07072__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__A top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold818 top.DUT.register\[16\]\[2\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_48_clk _00864_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 top.DUT.register\[1\]\[29\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_208_Right_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ clknet_leaf_43_clk _00795_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ _01898_ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__and2_1
XANTENNA__08887__B _03977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ _03849_ _03884_ net318 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XANTENNA__07780__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _02244_ _02638_ _02719_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__or3b_1
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07672_ top.DUT.register\[20\]\[10\] net560 net544 top.DUT.register\[24\]\[10\] _02788_
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a221o_1
XANTENNA__07532__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _04443_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06623_ _01713_ _01737_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ net131 _04370_ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_47_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06554_ top.DUT.register\[2\]\[0\] net684 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07312__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ net915 top.pc\[9\] net910 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07835__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06638__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06485_ _01388_ top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08224_ _03336_ _03339_ net317 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ _02153_ _03103_ _03157_ _03155_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__o31a_1
XFILLER_0_200_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07106_ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__inv_2
XANTENNA__09239__A _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07063__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ net829 _03202_ net468 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07037_ net298 _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06810__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout770_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _03371_ _01730_ _02880_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__mux2_1
XANTENNA__06598__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07939_ _02003_ _03053_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ net1468 net242 net481 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XANTENNA__06885__X _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ top.pc\[28\] _04606_ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_211_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10881_ net1422 net143 net492 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XANTENNA__06877__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12620_ clknet_leaf_3_clk _00166_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_195_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09815__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12551_ clknet_leaf_84_clk _00097_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[16\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11083__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _05352_ _05354_ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__a21o_2
X_12482_ clknet_leaf_90_clk _00029_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _05259_ _05261_ net478 _05231_ top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1
+ _05294_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__A1_N net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07054__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ _01393_ _01394_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10315_ net1664 net154 net521 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13103_ clknet_leaf_22_clk _00649_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11295_ net906 _05143_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_210_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ clknet_leaf_2_clk _00580_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ net163 top.DUT.register\[9\]\[25\] net385 vssd1 vssd1 vccd1 vccd1 _00403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net39 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
XANTENNA__09751__A1 _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ net1572 net161 net526 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06868__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ net1127 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13704__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12818_ clknet_leaf_106_clk _00364_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13798_ clknet_leaf_69_clk _01323_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ clknet_leaf_113_clk _00295_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06270_ net1382 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[28\] sky130_fd_sc_hd__and2_1
XANTENNA__07293__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08515__X _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__B2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold604 top.DUT.register\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold615 top.DUT.register\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold626 top.DUT.register\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold637 top.DUT.register\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold648 top.DUT.register\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_2
Xhold659 top.DUT.register\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _04942_ _04943_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_6_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11129__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _03007_ _03981_ _03008_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12641__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09891_ _04868_ _04873_ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10432__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ net473 _03927_ _03934_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07753__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08773_ _03330_ _03335_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout184_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07724_ _02839_ _02840_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__or2_2
XANTENNA__07505__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07655_ _02366_ _02769_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__or2_1
XANTENNA__06859__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08409__Y _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ net912 _01602_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07586_ top.DUT.register\[19\]\[15\] net673 net546 top.DUT.register\[24\]\[15\] _02702_
+ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a221o_1
XANTENNA__08138__A _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ net918 top.pc\[12\] _04367_ net911 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__o211a_1
X_06537_ net746 _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ net822 _04301_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_4_10__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ top.DUT.register\[6\]\[0\] net597 net593 top.DUT.register\[8\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a22o_1
XANTENNA__07284__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08481__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ _03321_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ _01411_ net853 _04224_ _04238_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__o22ai_1
XANTENNA__10607__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06399_ top.a1.instruction\[19\] net830 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__and2_1
X_08138_ _02195_ _03252_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout985_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08069_ top.DUT.register\[18\]\[17\] net660 net632 top.DUT.register\[27\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10100_ net201 net1321 net386 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XANTENNA__07992__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ net1165 net878 net846 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ net197 net2275 net530 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__09733__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10342__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11982_ _05819_ _05833_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_1
XANTENNA__07651__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ clknet_leaf_63_clk _01251_ net1106 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ net1834 net200 net485 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10864_ net1994 net213 net489 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__mux2_1
X_13652_ clknet_leaf_89_clk _01193_ net1013 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ clknet_leaf_0_clk _00149_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13583_ clknet_leaf_64_clk _01124_ net1097 vssd1 vssd1 vccd1 vccd1 top.a1.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10795_ net223 net2217 net410 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12534_ clknet_leaf_110_clk _00080_ net947 vssd1 vssd1 vccd1 vccd1 top.ramstore\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08472__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08472__B2 _03581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10517__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[28\] net1081 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[28\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07027__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _05264_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or2_2
X_12396_ net2253 net120 _00017_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11347_ net1247 net843 _05211_ net1115 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07983__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _05147_ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nor2_1
XANTENNA_output78_A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13017_ clknet_leaf_58_clk _00563_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10229_ net234 net1939 net384 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
XANTENNA__10252__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__B top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07127__A _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08160__B1 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ net305 net335 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ _02481_ _02483_ _02485_ _02487_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__or4_4
XANTENNA__06972__Y _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ _03961_ _04011_ _04056_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__and3_1
X_06322_ _01458_ _01332_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07266__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _03551_ _04092_ _04093_ _03468_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_40_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06253_ net1187 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[11\] sky130_fd_sc_hd__and2_1
XANTENNA__10427__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12838__RESET_B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07018__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06184_ top.lcd.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
Xhold401 top.DUT.register\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 top.DUT.register\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 top.DUT.register\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 top.DUT.register\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 top.DUT.register\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 top.DUT.register\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold467 top.DUT.register\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold478 top.DUT.register\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 top.DUT.register\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _04914_ _04916_ _04917_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12420__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
Xfanout925 _01400_ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_A _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_55_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10162__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout947 net949 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
X_09874_ _03879_ net455 net534 _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o211a_1
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_2
Xhold1101 top.DUT.register\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 net994 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 top.DUT.register\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08825_ net903 top.pc\[23\] net538 _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a22o_1
Xhold1123 top.DUT.register\[5\]\[9\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 top.DUT.register\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 top.DUT.register\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 top.DUT.register\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 top.DUT.register\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net277 _03852_ net271 _03681_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__o2bb2a_1
Xhold1178 top.DUT.register\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 top.ramload\[18\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
X_07707_ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__inv_2
X_08687_ net306 _03379_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06595__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07638_ top.DUT.register\[20\]\[8\] net562 net645 top.DUT.register\[10\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ _02679_ _02681_ _02683_ _02685_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ net915 top.pc\[11\] _04351_ net910 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__o211a_1
XANTENNA__07257__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ net158 net1625 net502 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07500__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06465__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _02448_ _02591_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__nand2_1
XANTENNA__10337__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ top.lcd.cnt_20ms\[5\] _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07009__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ top.a1.halfData\[5\] _01423_ _01427_ _01381_ _01420_ vssd1 vssd1 vccd1 vccd1
+ _05104_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_170_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12181_ _06037_ _06041_ _06040_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__a21boi_2
XANTENNA__09954__B2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net71 net881 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__and2_1
Xhold990 top.DUT.register\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ net9 net862 net834 net1348 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__o22a_1
XANTENNA__10072__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__B _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net242 net1880 net532 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
XANTENNA__13367__RESET_B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10800__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _05800_ _05801_ _05822_ _05824_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__a211o_1
XFILLER_0_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_74_clk _00016_ net1090 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_196_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _04181_ net617 _04958_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and3_4
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11896_ _05745_ _05746_ _05756_ _05754_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13635_ clknet_leaf_75_clk net1156 net1082 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net1388 _04941_ net493 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13566_ clknet_leaf_32_clk _01112_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ net158 net1804 net371 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06456__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ clknet_leaf_92_clk _00063_ net997 vssd1 vssd1 vccd1 vccd1 top.ramstore\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10247__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ clknet_leaf_58_clk _01043_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12448_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[11\] net1077 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[11\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09945__A1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12379_ top.pad.button_control.r_counter\[13\] _06153_ vssd1 vssd1 vccd1 vccd1 _06155_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09337__A _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07420__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ top.DUT.register\[10\]\[22\] net727 net759 top.DUT.register\[2\]\[22\] _02056_
+ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09771__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ top.DUT.register\[21\]\[25\] net611 net763 top.DUT.register\[30\]\[25\] _01987_
+ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a221o_1
XFILLER_0_206_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08610_ net467 _03713_ _03711_ _03709_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_128_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ net132 _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08541_ net1359 net858 net836 _03647_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ net904 top.pc\[7\] net538 _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07423_ top.DUT.register\[22\]\[5\] net555 net665 top.DUT.register\[14\]\[5\] _02539_
+ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a221o_1
XANTENNA__06695__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_A _04941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ top.DUT.register\[12\]\[5\] net737 net710 top.DUT.register\[7\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a22o_1
XANTENNA__12232__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08416__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06305_ net1238 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[31\] sky130_fd_sc_hd__and2_1
XFILLER_0_33_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10157__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ top.DUT.register\[26\]\[2\] net721 net717 top.DUT.register\[9\]\[2\] _02401_
+ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout314_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ _03051_ _04083_ net1630 net891 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06236_ top.Ren top.Wen vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 top.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A1 _03995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06167_ top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold231 top.DUT.register\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold242 top.DUT.register\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 top.DUT.register\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07947__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 top.DUT.register\[13\]\[8\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold275 top.DUT.register\[16\]\[22\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout683_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold286 top.DUT.register\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _01660_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_4
Xhold297 top.a1.row2\[1\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
X_09926_ net160 net2182 net392 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
Xfanout722 _01548_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_2
Xfanout733 _01540_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 _04726_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_2
Xfanout755 _01575_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
Xfanout766 _01560_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
XANTENNA_fanout850_A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 _01555_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
X_09857_ net190 net1447 net390 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__mux2_1
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 _01644_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_2
X_08808_ net279 net356 vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__or2_1
XANTENNA__10620__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ top.pc\[13\] _04378_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ _03158_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_1_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _05562_ _05574_ _05607_ _05609_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__or4_1
XANTENNA__07478__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ net1371 net204 net499 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11681_ net178 _05537_ _05538_ _05504_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ clknet_leaf_2_clk _00966_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ net217 net1980 net374 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XANTENNA__12223__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07230__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ net230 net2251 net503 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__mux2_1
X_13351_ clknet_leaf_52_clk _00897_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ top.lcd.cnt_500hz\[0\] net742 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10494_ net246 net1473 net380 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
X_13282_ clknet_leaf_11_clk _00828_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12233_ net1107 _04674_ net870 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12164_ _06009_ _06020_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09157__A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net923 net1337 net875 _05057_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ _05940_ _05941_ _05930_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a21o_1
XANTENNA_input32_X net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11046_ top.busy_o net852 wb.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_207_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10530__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12997_ clknet_leaf_40_clk _00543_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ _05776_ _05784_ _05796_ _05797_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__and4_1
XFILLER_0_157_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06677__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11879_ _01398_ net127 vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ clknet_leaf_93_clk _01159_ net996 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13549_ clknet_leaf_114_clk _01095_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07070_ _02180_ _02182_ _02184_ _02186_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__or4_1
XANTENNA__09148__C_N _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07641__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10705__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07929__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07972_ top.DUT.register\[3\]\[18\] net691 net643 top.DUT.register\[10\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ top.pc\[1\] _04721_ _04723_ _04725_ net911 vssd1 vssd1 vccd1 vccd1 _00121_
+ sky130_fd_sc_hd__o221a_1
X_06923_ top.DUT.register\[28\]\[23\] net738 net766 top.DUT.register\[11\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
XANTENNA__10440__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ _01417_ _04656_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__xnor2_1
X_06854_ _01964_ _01966_ _01968_ _01970_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__or4_1
X_06785_ top.DUT.register\[30\]\[30\] net763 net714 top.DUT.register\[25\]\[30\] _01901_
+ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a221o_1
X_09573_ top.pc\[26\] _04576_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o21ai_2
XANTENNA__08106__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_A _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _03400_ _03570_ _03628_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__o21a_1
XANTENNA__08657__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08657__B2 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06668__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _03450_ _03562_ net290 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout431_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _02517_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08386_ _03302_ _03340_ net288 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08409__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ top.DUT.register\[26\]\[6\] net721 net772 top.DUT.register\[27\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07093__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ _02378_ _02380_ _02382_ _02384_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__or4_1
XANTENNA__07632__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06219_ _00009_ top.a1.nextHex\[7\] vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[2\] sky130_fd_sc_hd__or2_1
X_09007_ _02767_ net620 net1372 net887 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06840__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ top.DUT.register\[12\]\[10\] net734 net592 top.DUT.register\[8\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XANTENNA__10615__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07396__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 net532 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_8
Xfanout541 _01692_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_8
Xfanout552 net553 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_4
X_09909_ top.pc\[25\] _04576_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and2_1
Xfanout563 _01673_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_2
Xfanout574 _01657_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net587 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_8
X_12920_ clknet_leaf_36_clk _00466_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_4
XANTENNA__10350__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__B _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07699__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ clknet_leaf_110_clk _00397_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_202_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _05650_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12782_ clknet_leaf_96_clk _00328_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09845__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11733_ _05586_ _05590_ _05593_ _05584_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12523__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11664_ _05486_ _05524_ _05523_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_126_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13403_ clknet_leaf_1_clk _00949_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ net150 net2128 net423 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ _05443_ _05448_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__a21o_1
XANTENNA__07084__A0 _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ clknet_leaf_104_clk _00880_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10546_ net163 net2281 net429 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__mux2_1
XANTENNA__07623__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06831__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13265_ clknet_leaf_10_clk _00811_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10525__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10477_ net175 net1414 net506 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13650__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ net1440 net866 net831 _06021_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13196_ clknet_leaf_4_clk _00742_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08997__Y _04082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12147_ top.a1.dataIn\[3\] _05981_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__nand2_1
XANTENNA__09615__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ _05909_ _05916_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09533__C1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ top.a1.dataIn\[8\] net869 net864 _05041_ vssd1 vssd1 vccd1 vccd1 _05042_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06898__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06570_ _01650_ _01676_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__nor2_4
XANTENNA__09836__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08240_ _03341_ _03355_ net302 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08171_ _01720_ _01727_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07122_ top.DUT.register\[21\]\[14\] net609 net770 top.DUT.register\[27\]\[14\] _02238_
+ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07075__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ top.DUT.register\[21\]\[17\] net609 net751 top.DUT.register\[19\]\[17\] _02169_
+ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10435__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__Y _03800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ top.DUT.register\[11\]\[20\] net700 net692 top.DUT.register\[3\]\[20\] _03071_
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_182_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06906_ _02013_ _02022_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__nor2_8
XANTENNA__10170__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ net825 _03002_ _02617_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06889__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ top.pc\[30\] _04638_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__or2_1
X_06837_ top.DUT.register\[14\]\[27\] net792 net760 top.DUT.register\[30\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout646_A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _04583_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__or2_1
X_06768_ top.DUT.register\[25\]\[29\] net711 net758 top.DUT.register\[2\]\[29\] _01884_
+ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10437__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ top.pc\[22\] _04511_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06699_ top.DUT.register\[7\]\[4\] net574 net673 top.DUT.register\[19\]\[4\] _01815_
+ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08438_ net904 top.pc\[6\] net537 _03548_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a22o_1
XANTENNA__07853__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08369_ net469 _02518_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07066__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ net1501 net217 net513 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09259__X _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _05240_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__inv_2
XANTENNA__08802__A1 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ net1821 net228 net519 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__mux2_1
XANTENNA__10345__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10262_ net238 net2159 net436 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__mux2_1
X_13050_ clknet_leaf_20_clk _00596_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ _05837_ _05841_ _05858_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__and3_1
XANTENNA__08030__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ net244 net2296 net440 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
XFILLER_0_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout371 _04997_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10080__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 _04978_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_6
Xfanout393 _04734_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12903_ clknet_leaf_49_clk _00449_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12834_ clknet_leaf_25_clk _00380_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09441__Y _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12765_ clknet_leaf_118_clk _00311_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08097__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11716_ _05571_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__and2_1
XANTENNA__07844__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ clknet_leaf_33_clk _00242_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ _05497_ _05498_ _05507_ _05488_ _05480_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a2111o_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XFILLER_0_140_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11578_ _05401_ _05435_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__xor2_1
X_13317_ clknet_leaf_40_clk _00863_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold808 top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10255__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__B _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10529_ net235 net1567 net428 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__mux2_1
Xhold819 top.DUT.register\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12036__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13248_ clknet_leaf_105_clk _00794_ net981 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08021__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ clknet_leaf_5_clk _00725_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06583__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _02664_ _02855_ _02856_ _02825_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07671_ top.DUT.register\[1\]\[10\] net703 net627 top.DUT.register\[29\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a22o_1
X_09410_ _02174_ _04445_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__xnor2_1
X_06622_ net366 net297 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__and2_1
XANTENNA__12445__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09341_ net135 _04375_ _04382_ net821 net915 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o221a_1
X_06553_ net746 _01647_ _01652_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__and3_4
XPHY_EDGE_ROW_188_Left_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07296__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__B _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06991__X _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ net131 _04310_ net915 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06484_ _01388_ top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07835__A2 _02951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08223_ _03337_ _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout227_A _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _03079_ _03131_ _02109_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07105_ _02212_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__nor2_4
XFILLER_0_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10165__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ _03192_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__nor2_4
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07036_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout596_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09526__Y _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__Y _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ net473 _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_149_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07938_ _02003_ _03052_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07869_ top.DUT.register\[14\]\[27\] net663 net647 top.DUT.register\[12\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ top.pc\[28\] _04606_ _04618_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a21o_1
X_10880_ net1854 net148 net489 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09539_ top.pc\[25\] _04557_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nor2_1
XANTENNA__08079__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ clknet_leaf_84_clk _00096_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07287__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _05358_ _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__nand2_1
X_12481_ clknet_leaf_90_clk _00028_ net1010 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07039__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _05265_ _05278_ _05283_ _05286_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__o41ai_4
XTAP_TAPCELL_ROW_78_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10075__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ top.a1.dataIn\[18\] top.a1.dataIn\[19\] top.a1.dataIn\[17\] top.a1.dataIn\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13102_ clknet_leaf_96_clk _00648_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ net1768 net160 net523 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11294_ net1174 net844 _05164_ net1115 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_210_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ clknet_leaf_28_clk _00579_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10245_ net168 net1495 net384 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XANTENNA__10803__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08003__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1104 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1111 net1121 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_2
XANTENNA__07211__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net2163 net162 net528 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09751__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_201_Left_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout190 _04851_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09171__Y _04224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08509__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12817_ clknet_leaf_9_clk _00363_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13797_ clknet_leaf_69_clk _01322_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07278__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ clknet_leaf_3_clk _00294_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07817__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_210_Left_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ clknet_leaf_56_clk _00225_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08244__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold605 top.DUT.register\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold616 top.DUT.register\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 top.DUT.register\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 top.DUT.register\[8\]\[22\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold649 top.DUT.register\[17\]\[13\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08910_ net1283 net861 net838 _03999_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a22o_1
XANTENNA__09727__C1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10713__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ top.pc\[23\] _02615_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07202__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ _03032_ net459 _03929_ _02523_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a221o_1
XANTENNA__09742__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13593__Q top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ net307 _03504_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07723_ _02489_ _02549_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout177_A _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07654_ _02366_ _02768_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06605_ _01387_ _01603_ _01716_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__or3b_1
X_07585_ top.DUT.register\[13\]\[15\] net677 net653 top.DUT.register\[17\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11065__A1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ net133 _04352_ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06536_ top.a1.instruction\[21\] net799 top.a1.instruction\[20\] vssd1 vssd1 vccd1
+ vccd1 _01653_ sky130_fd_sc_hd__and3b_2
XFILLER_0_8_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ _04286_ _04289_ _04300_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ _01574_ _01577_ _01580_ _01583_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__or4_1
XFILLER_0_211_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ net323 _02469_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_190_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ net138 _04227_ _04228_ _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__o31a_1
X_06398_ _01485_ _01514_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ net352 _03252_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08068_ top.DUT.register\[8\]\[17\] net557 net628 top.DUT.register\[29\]\[17\] _03184_
+ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06795__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ top.DUT.register\[28\]\[18\] net738 net784 top.DUT.register\[29\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
XANTENNA__10623__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ net201 net2260 net529 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06402__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09713__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _05819_ _05833_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13720_ clknet_leaf_63_clk _01250_ net1106 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10932_ net1477 net203 net487 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ clknet_leaf_110_clk net1224 net947 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
X_10863_ net1593 net217 net489 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11056__A1 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ clknet_leaf_15_clk _00148_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ clknet_leaf_64_clk _01123_ net1097 vssd1 vssd1 vccd1 vccd1 top.a1.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ net229 net1613 net412 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07520__X _02637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__C _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12533_ clknet_leaf_89_clk _00079_ net1016 vssd1 vssd1 vccd1 vccd1 top.ramstore\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12464_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[27\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08064__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13678__Q net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ _05246_ net478 _05236_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10567__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ net2309 net119 _00017_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ top.a1.row1\[60\] _05140_ _05210_ net845 vssd1 vssd1 vccd1 vccd1 _05211_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08351__X _03465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06786__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10533__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ top.lcd.nextState\[5\] top.lcd.nextState\[4\] _05137_ vssd1 vssd1 vccd1 vccd1
+ _05148_ sky130_fd_sc_hd__or3_1
XANTENNA__09185__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ clknet_leaf_37_clk _00562_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ net238 net1991 net385 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07735__A1 _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06538__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 top.pad.button_control.debounce vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net1901 net233 net527 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ clknet_leaf_59_clk _01372_ net1102 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09061__C _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11047__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07370_ top.DUT.register\[22\]\[5\] net606 net775 top.DUT.register\[2\]\[5\] _02486_
+ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06321_ net901 net845 net844 top.lcd.currentState\[2\] net1114 vssd1 vssd1 vccd1
+ vccd1 _01332_ sky130_fd_sc_hd__o221a_2
XFILLER_0_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10708__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09040_ _03497_ _03524_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nand2_1
X_06252_ net2232 net894 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[10\] sky130_fd_sc_hd__and2_1
XANTENNA__07671__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06183_ top.pad.button_control.r_counter\[8\] vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_107_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09412__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09412__B2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 top.DUT.register\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 top.DUT.register\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07423__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 top.DUT.register\[11\]\[29\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 top.DUT.register\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 top.DUT.register\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06777__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 top.DUT.register\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 top.DUT.register\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold479 top.DUT.register\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10443__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
Xfanout915 net917 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
Xfanout926 net928 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 net942 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_2
X_09873_ _04862_ _04863_ _04864_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a211o_1
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout959 net960 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_2
X_08824_ _03367_ _03900_ _03912_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__a211o_1
Xhold1102 top.DUT.register\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07037__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1113 top.DUT.register\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 top.DUT.register\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 top.DUT.register\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 top.DUT.register\[20\]\[10\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _03769_ _03851_ net290 vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_116_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1157 top.DUT.register\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1179 top.DUT.register\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07706_ _02821_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_179_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ net304 _03356_ _03571_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07637_ top.DUT.register\[6\]\[8\] net578 _02753_ vssd1 vssd1 vccd1 vccd1 _02754_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07988__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ top.DUT.register\[4\]\[9\] net550 net625 top.DUT.register\[16\]\[9\] _02684_
+ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ net135 _04341_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__o21ai_1
X_06519_ top.a1.instruction\[8\] _01486_ net824 top.a1.instruction\[13\] vssd1 vssd1
+ vccd1 vccd1 _01636_ sky130_fd_sc_hd__a22o_1
XANTENNA__10618__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ net857 _01752_ _02614_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_118_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07662__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ _02448_ _02591_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_125_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09169_ _01410_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11200_ top.a1.row1\[61\] _05096_ _05103_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__o21a_1
XANTENNA__07414__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12180_ _06023_ _06038_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06768__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ net924 net1306 net876 _05065_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a31o_1
XANTENNA__10353__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 top.DUT.register\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 top.DUT.register\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ net8 net862 net834 net1429 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__o22a_1
X_10013_ net615 _04962_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_134_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07193__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06940__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _05822_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__or2_1
X_13703_ clknet_leaf_74_clk _00015_ net1089 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10915_ net1637 net139 net408 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
X_11895_ _05690_ _05714_ _05727_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11029__A1 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12226__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ clknet_leaf_91_clk _01175_ net1003 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
X_10846_ net1350 net150 net495 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13565_ clknet_leaf_1_clk _01111_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_Left_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10777_ net165 net1689 net373 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10528__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12516_ clknet_leaf_93_clk _00062_ net995 vssd1 vssd1 vccd1 vccd1 top.ramstore\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13496_ clknet_leaf_36_clk _01042_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12447_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[10\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09618__A _01898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ _06153_ _06154_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06759__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ top.a1.row1\[3\] _05154_ _05158_ top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1
+ _05197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10263__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09337__B _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09905__X _04895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ top.DUT.register\[14\]\[25\] net795 net782 top.DUT.register\[3\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08381__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ net902 top.pc\[10\] net537 _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ net463 _03551_ _03575_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a211o_2
XFILLER_0_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07422_ top.DUT.register\[30\]\[5\] net698 net563 top.DUT.register\[20\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13077__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09800__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07601__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07353_ net321 _02468_ _02449_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10438__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06304_ net1524 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[30\] sky130_fd_sc_hd__and2_1
XANTENNA__07644__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07284_ top.DUT.register\[28\]\[2\] net740 net786 top.DUT.register\[29\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06998__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09023_ _03028_ net621 net1328 net891 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a2bb2o_1
X_06235_ net1 net877 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout307_A _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1__f_clk_X clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 top.DUT.register\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09528__A _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 top.DUT.register\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06166_ net912 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold232 top.DUT.register\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold265 top.DUT.register\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 top.DUT.register\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08151__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 top.DUT.register\[27\]\[9\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout701 _01660_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09815__X _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout712 _01567_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
X_09925_ _03977_ net456 net536 _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o211a_2
Xhold298 top.DUT.register\[1\]\[28\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout723 _01546_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_8
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
XANTENNA__11793__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout676_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _04726_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_1
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
X_09856_ _03838_ net454 net533 _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__o211a_2
Xfanout767 _01560_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
XANTENNA__10901__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06887__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 net791 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
X_08807_ _03557_ _03558_ net310 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__o21a_1
XANTENNA__09263__A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ net218 net2053 net391 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ top.DUT.register\[29\]\[19\] net784 _02114_ _02115_ vssd1 vssd1 vccd1 vccd1
+ _02116_ sky130_fd_sc_hd__a211o_1
XANTENNA__06922__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _03105_ _03806_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nand2_1
XANTENNA__09004__A1_N _02548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08669_ _03680_ _03768_ net289 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09872__A1 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ net1236 net210 net497 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06686__A1 top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ _05518_ _05536_ _05539_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__and3_1
XANTENNA__07883__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09019__A1_N net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ net222 net1504 net375 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10348__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13350_ clknet_leaf_47_clk _00896_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07230__B _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10562_ net234 net2070 net503 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12301_ net1119 _01453_ _06080_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11968__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ clknet_leaf_42_clk _00827_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10493_ net249 net1907 net380 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
X_12232_ net1356 net868 net833 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__a21o_1
XANTENNA__09927__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12163_ _06009_ _06020_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__or2_1
XANTENNA__09157__B _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07229__Y _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ net40 net882 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and2_1
XANTENNA__09725__X _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ _05936_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_207_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ top.busy_o wb.prev_BUSY_O net863 vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_207_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10811__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08363__A1 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06913__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__B _01733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12996_ clknet_leaf_28_clk _00542_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_clk_X clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _05777_ _05783_ _05795_ _05798_ _05780_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_28_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08666__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A1 _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07874__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _05701_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__xnor2_2
X_13617_ clknet_leaf_74_clk _01158_ net1087 vssd1 vssd1 vccd1 vccd1 top.ramload\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10258__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829_ net1400 net221 net494 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09076__C1 _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08236__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13548_ clknet_leaf_2_clk _01094_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_49_clk _01025_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09379__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08252__A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08051__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _03085_ _03086_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_52_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ _04085_ _04724_ _04721_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__a21bo_1
X_06922_ top.DUT.register\[4\]\[23\] net580 net758 top.DUT.register\[2\]\[23\] _02038_
+ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a221o_1
XANTENNA__10721__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ top.pc\[30\] _04643_ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__o21a_1
X_06853_ top.DUT.register\[22\]\[26\] net606 net780 top.DUT.register\[1\]\[26\] _01969_
+ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a221o_1
XANTENNA__09712__C_N _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ top.pc\[26\] _04576_ _04586_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a21o_1
X_06784_ top.DUT.register\[27\]\[30\] net773 net710 top.DUT.register\[7\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08523_ _03617_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11110__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__A1 _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _03449_ _03563_ net290 vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07405_ _01719_ _01733_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__or2_4
XANTENNA__07331__A _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08385_ _02841_ _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10168__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09957__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07336_ top.DUT.register\[20\]\[6\] net591 net710 top.DUT.register\[7\]\[6\] _02452_
+ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a221o_1
XANTENNA__07617__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08290__A0 _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07267_ top.DUT.register\[20\]\[3\] net590 net757 top.DUT.register\[3\]\[3\] _02383_
+ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ _02610_ net621 net1227 net890 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__a2bb2o_1
X_06218_ _01433_ top.a1.hexop\[4\] _01428_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[1\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06234__X _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07198_ top.DUT.register\[21\]\[10\] net608 net754 top.DUT.register\[18\]\[10\] _02314_
+ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout793_A _01529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__B2 _02284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout960_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _04983_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_6
Xfanout542 _01692_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10631__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ top.pc\[24\] _04557_ _04892_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a21oi_1
Xfanout553 net555 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_4
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_8
Xfanout575 _01657_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_8
X_09839_ net819 _04453_ _04834_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__o21ba_1
Xfanout597 net599 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_4
XFILLER_0_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ clknet_leaf_105_clk _00396_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13610__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11801_ _05629_ net130 _05620_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_202_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ clknet_leaf_115_clk _00327_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09845__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ _05553_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07856__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A _01775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11663_ _05483_ _05505_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10078__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13402_ clknet_leaf_14_clk _00948_ net987 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10614_ net156 net2009 net423 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
Xwire921 _01419_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09073__A2 _03541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11594_ _05425_ _05450_ _05453_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_141_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ clknet_leaf_101_clk _00879_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ net166 net1700 net429 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__mux2_1
XANTENNA__10806__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ clknet_leaf_117_clk _00810_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10476_ net179 net1711 net506 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__mux2_1
XANTENNA__13686__Q top.pc\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12306__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net1891 net867 net831 _06032_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ clknet_leaf_4_clk _00741_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07387__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _05999_ _06006_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10541__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _05918_ _05935_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07139__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ top.a1.data\[4\] top.a1.dataInTemp\[8\] net796 vssd1 vssd1 vccd1 vccd1 _05041_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12979_ clknet_leaf_108_clk _00525_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09836__A1 _03800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08170_ _01941_ _02878_ _03268_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07121_ top.DUT.register\[18\]\[14\] net779 net761 top.DUT.register\[30\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08811__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07052_ top.DUT.register\[29\]\[17\] net785 net713 top.DUT.register\[25\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__clkbuf_4
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07378__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09772__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10451__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ top.DUT.register\[17\]\[20\] net652 net644 top.DUT.register\[10\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_182_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06905_ _02017_ _02019_ _02021_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__or3_2
XFILLER_0_128_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07885_ _02992_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__or2_4
XFILLER_0_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06230__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ top.pc\[30\] _04638_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nand2_1
X_06836_ _01946_ _01948_ _01950_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__or4_1
XFILLER_0_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09555_ top.pc\[26\] _04565_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__nor2_1
X_06767_ top.DUT.register\[28\]\[29\] net738 net760 top.DUT.register\[30\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout541_A _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout639_A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net303 _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or2_1
XANTENNA__09260__B _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09486_ _04506_ _04507_ _04505_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06698_ top.DUT.register\[1\]\[4\] net705 net685 top.DUT.register\[2\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a22o_1
XANTENNA__07302__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ net462 _03524_ _03547_ net464 _03544_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08368_ net271 _03478_ _03479_ _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o22a_1
XFILLER_0_190_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07319_ top.DUT.register\[2\]\[7\] net774 net764 top.DUT.register\[19\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08299_ net292 _03412_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__nand2_1
XANTENNA__12213__A2_N _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ net1617 net233 net519 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ net245 net1958 net436 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__mux2_1
X_12000_ _05826_ _05835_ _05836_ _05825_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07369__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11165__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ net249 net1936 net440 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
XANTENNA__06577__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10361__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__B _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_1
XANTENNA__13109__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 _04997_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_8
Xfanout383 _04978_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_4
Xfanout394 _02521_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
X_12902_ clknet_leaf_48_clk _00448_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ clknet_leaf_49_clk _00379_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11045__X _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07829__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ clknet_leaf_51_clk _00310_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _05574_ _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ clknet_leaf_112_clk _00241_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11646_ _05453_ _05484_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_1
XFILLER_0_181_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
Xinput36 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_103_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10536__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ top.a1.dataIn\[13\] _05435_ _05436_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13316_ clknet_leaf_28_clk _00862_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10528_ net236 net1692 net428 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__mux2_1
Xhold809 top.DUT.register\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_47_clk _00793_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08006__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__C1 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ net254 net1852 net507 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__mux2_1
XANTENNA__08557__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ clknet_leaf_14_clk _00724_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06568__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _05952_ _05986_ _05951_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10271__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__B _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ top.DUT.register\[17\]\[10\] net651 net643 top.DUT.register\[10\]\[10\] _02786_
+ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a221o_1
XFILLER_0_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07532__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07433__X _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ net366 net297 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__or2_1
XANTENNA__08248__Y _03364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ _04376_ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06552_ net747 _01649_ _01656_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ net135 _04309_ _04316_ net821 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__o22a_1
X_06483_ net914 net913 _01484_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__and3_2
XFILLER_0_173_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ net325 _02153_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12414__RESET_B net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ _02881_ _02902_ _03269_ _02878_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10446__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07104_ _02214_ _02216_ _02218_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__or4_2
XANTENNA__08796__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _03194_ _03196_ _03198_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or4_2
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ _02150_ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout1031_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09095__X _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09745__B1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net306 _03752_ _03908_ net269 _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_149_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07771__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__X _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06598__C top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _02003_ _03052_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__and2_2
XFILLER_0_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ top.DUT.register\[9\]\[27\] net639 net627 top.DUT.register\[29\]\[27\] _02984_
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ _04631_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__nand2_1
X_06819_ top.DUT.register\[26\]\[31\] net722 net718 top.DUT.register\[9\]\[31\] _01935_
+ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a221o_1
XANTENNA__06731__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ top.DUT.register\[4\]\[29\] net548 net651 top.DUT.register\[17\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09538_ net134 _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09469_ top.pc\[21\] _04484_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11083__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11500_ _05359_ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ clknet_leaf_89_clk _00027_ net1015 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ _05289_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10356__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12137__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11362_ top.a1.dataIn\[31\] top.a1.dataIn\[30\] _05222_ vssd1 vssd1 vccd1 vccd1 _05223_
+ sky130_fd_sc_hd__nand3_1
XANTENNA__06798__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ clknet_leaf_113_clk _00647_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10313_ net1790 net162 net524 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ top.a1.row1\[120\] _05129_ _05135_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_91_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_210_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13032_ clknet_leaf_31_clk _00578_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10244_ net173 net2237 net382 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
Xfanout1101 net1104 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ net2164 net167 net527 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
Xfanout180 _04867_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_1
XANTENNA__06970__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 _04841_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07514__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ net1126 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
X_12816_ clknet_leaf_117_clk _00362_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13796_ clknet_leaf_69_clk _01321_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12747_ clknet_leaf_4_clk _00293_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ clknet_leaf_19_clk _00224_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08525__A _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11629_ _05456_ _05465_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10266__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08778__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__B2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold606 top.DUT.register\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold617 top.DUT.register\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 top.DUT.register\[17\]\[31\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
XANTENNA_max_cap342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 top.DUT.register\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11129__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__Y _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ net276 _01941_ net395 _03030_ net477 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_29_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07753__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ _03132_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08950__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06961__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _02489_ _02549_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07505__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__B2 _03801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _02366_ _02768_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__nor2_1
X_06604_ _01607_ _01717_ _01599_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07584_ top.DUT.register\[11\]\[15\] net701 _02700_ vssd1 vssd1 vccd1 vccd1 _02701_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09258__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ net137 _04357_ _04365_ net822 net918 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__o221a_1
X_06535_ top.a1.instruction\[22\] top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_38_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _04286_ _04289_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06466_ top.DUT.register\[13\]\[0\] net789 net716 top.DUT.register\[9\]\[0\] _01582_
+ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ net322 _02489_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ net823 _04235_ _04236_ net134 _04231_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__o32a_1
X_06397_ _01482_ _01512_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_190_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ net352 _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__nor2_1
XANTENNA__09966__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08067_ top.DUT.register\[6\]\[17\] net577 net624 top.DUT.register\[16\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__a22o_1
XANTENNA__10904__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ top.DUT.register\[1\]\[18\] net781 net707 top.DUT.register\[7\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
XANTENNA__09266__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A _04224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07057__Y _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06436__A_N top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07744__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A1_N net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _02927_ _02954_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _05812_ _05839_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_197_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08169__X _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net2140 net208 net485 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
XANTENNA__06704__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10862_ top.DUT.register\[28\]\[11\] net219 net490 vssd1 vssd1 vccd1 vccd1 _00997_
+ sky130_fd_sc_hd__mux2_1
X_13650_ clknet_leaf_75_clk net1163 net1083 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ clknet_leaf_59_clk _00147_ net1103 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ clknet_leaf_64_clk _01122_ net1097 vssd1 vssd1 vccd1 vccd1 top.a1.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ net232 net2030 net412 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12532_ clknet_leaf_93_clk _00078_ net995 vssd1 vssd1 vccd1 vccd1 top.ramstore\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06417__X _01534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08345__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10086__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ clknet_leaf_74_clk top.ru.next_FetchedInstr\[26\] net1088 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08064__B _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ _05238_ _05266_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__xor2_4
XFILLER_0_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09728__X _04742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ net2222 net118 _00017_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11345_ _05127_ _05153_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__nor2_1
XANTENNA__07432__A1 _02548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07983__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ net906 net900 vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__nand2_1
X_13015_ clknet_leaf_114_clk _00561_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ net244 net1641 net384 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ net1499 net238 net527 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 top.lcd.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06943__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10089_ net251 top.DUT.register\[5\]\[5\] net388 vssd1 vssd1 vccd1 vccd1 _00255_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06739__S net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13848_ clknet_leaf_59_clk _01371_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13066__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ clknet_leaf_64_clk _01304_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_06320_ top.lcd.nextState\[1\] _01453_ net844 net2219 net1118 vssd1 vssd1 vccd1 vccd1
+ _01331_ sky130_fd_sc_hd__o221a_2
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08255__A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06251_ net1653 net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[9\] sky130_fd_sc_hd__and2_1
XFILLER_0_143_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__C1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06182_ net1151 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold403 top.DUT.register\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 top.DUT.register\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10724__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 top.DUT.register\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 top.DUT.register\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold447 top.DUT.register\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold458 top.DUT.register\[5\]\[12\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 top.DUT.register\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ top.pc\[28\] _04622_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout905 top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _04511_ net361 net328 top.a1.dataIn\[21\] net363 vssd1 vssd1 vccd1 vccd1
+ _04865_ sky130_fd_sc_hd__a221o_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
Xhold1103 top.DUT.register\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ net465 _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_146_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 top.pad.keyCode\[7\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1125 top.DUT.register\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 top.DUT.register\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net316 _03809_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o21ai_1
Xhold1147 top.DUT.register\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 top.DUT.register\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 top.pad.button_control.r_counter\[7\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ net349 _02820_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08685_ _03208_ _03783_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_179_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_92_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ top.DUT.register\[8\]\[8\] net558 net546 top.DUT.register\[24\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_192_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08439__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ top.DUT.register\[6\]\[9\] net578 net665 top.DUT.register\[14\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_192_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_A _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout719_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ net131 _04336_ _04348_ _04349_ net915 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__o221a_1
X_06518_ net912 net824 _01634_ top.a1.instruction\[20\] _01631_ vssd1 vssd1 vccd1
+ vccd1 _01635_ sky130_fd_sc_hd__a221o_2
XANTENNA__07111__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07498_ _01613_ _01752_ _02614_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__o21a_2
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _02469_ _02567_ _04273_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06465__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06449_ net811 _01562_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_157_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ _04219_ _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__nand2_1
X_08119_ top.DUT.register\[7\]\[16\] net572 net564 top.DUT.register\[23\]\[16\] _03235_
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09099_ _02639_ _02663_ _02691_ _02716_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__and4_1
XANTENNA__10634__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11130_ net70 net882 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__and2_1
Xhold970 top.DUT.register\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 top.DUT.register\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ net7 net851 net850 top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__a22o_1
Xhold992 top.DUT.register\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07178__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ top.a1.instruction\[9\] top.a1.instruction\[10\] _04183_ net744 vssd1 vssd1
+ vccd1 vccd1 _04962_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_110_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09443__B _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11963_ _05787_ _05798_ _05793_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_83_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13702_ clknet_leaf_74_clk _00014_ net1089 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10914_ net1387 net145 net408 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11894_ _05690_ _05727_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12226__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13633_ clknet_leaf_111_clk net1217 net947 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10845_ net1797 net155 net493 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XANTENNA__10809__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10776_ net166 net1699 net373 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
X_13564_ clknet_leaf_19_clk _01110_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07102__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ clknet_leaf_93_clk _00061_ net996 vssd1 vssd1 vccd1 vccd1 top.ramstore\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06456__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ clknet_leaf_107_clk _01041_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[9\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12377_ net1332 _06151_ net815 vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10544__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09618__B _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ top.a1.row2\[43\] _05157_ _05165_ top.lcd.nextState\[0\] _05195_ vssd1 vssd1
+ vccd1 vccd1 _05196_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11259_ net906 top.lcd.nextState\[4\] top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1
+ _05130_ sky130_fd_sc_hd__and3b_1
XANTENNA__08905__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06916__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08470_ net464 _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_141_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07421_ _02531_ _02533_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06695__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10719__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07352_ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06303_ net1196 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[29\] sky130_fd_sc_hd__and2_1
X_07283_ top.DUT.register\[22\]\[2\] net605 net723 top.DUT.register\[16\]\[2\] _02399_
+ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ net1291 net888 _03177_ net622 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06234_ wb.curr_state\[1\] wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__or2_2
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold200 top.DUT.register\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold211 top.DUT.register\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ net911 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout202_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 top.a1.hexop\[1\] vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 top.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07947__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 top.DUT.register\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 top.DUT.register\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 top.DUT.register\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 top.DUT.register\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 top.DUT.register\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold299 top.DUT.register\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _04908_ _04909_ _04911_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o21ai_1
Xfanout702 _01660_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_4
Xfanout713 _01567_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1111_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_8
Xfanout735 net737 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_8
Xfanout746 _01646_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_2
XANTENNA__09544__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ net816 _04847_ _04848_ _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a211o_1
Xfanout757 _01570_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout571_A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _01560_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06887__B _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 _01541_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout669_A _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _03183_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__xnor2_1
X_06998_ top.DUT.register\[28\]\[19\] net738 net734 top.DUT.register\[12\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
X_09786_ _03695_ net454 net533 _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__o211a_2
XANTENNA__07580__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ net473 _03828_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_65_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07619_ top.DUT.register\[15\]\[11\] net688 net640 top.DUT.register\[9\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ net284 _03701_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ net224 net2271 net374 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10561_ net239 net1806 net504 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net1142 _06105_ _06106_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_20_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13280_ clknet_leaf_13_clk _00826_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10492_ net254 net1645 net380 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ top.a1.row2\[15\] net870 _05094_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__o21a_1
XANTENNA__10364__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06414__Y _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12162_ _05997_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__xnor2_2
X_11113_ net1223 net878 net846 top.ramstore\[31\] vssd1 vssd1 vccd1 vccd1 _01192_
+ sky130_fd_sc_hd__a22o_1
X_12093_ _05918_ _05935_ _05909_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ net1 wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_207_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__A1 top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09741__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ clknet_leaf_35_clk _00541_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_56_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09901__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946_ _05777_ _05795_ _05798_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12559__SET_B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06677__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10539__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _05700_ net127 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13616_ clknet_leaf_74_clk _01157_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramload\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ net2317 net223 net493 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ clknet_leaf_4_clk _01093_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ net236 net2133 net372 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XANTENNA__13104__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13478_ clknet_leaf_21_clk _01024_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10274__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12429_ clknet_leaf_78_clk top.ru.next_FetchedData\[24\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[24\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07929__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09916__X _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ top.DUT.register\[7\]\[18\] net572 net651 top.DUT.register\[17\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06921_ top.DUT.register\[12\]\[23\] net734 net711 top.DUT.register\[25\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__B1 _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_06852_ top.DUT.register\[5\]\[26\] net602 net728 top.DUT.register\[10\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
X_09640_ top.pc\[30\] _04643_ _04652_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a21o_1
XANTENNA__07562__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ _04597_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__nand2_1
X_06783_ net319 _01879_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08106__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ _03404_ _03570_ _03628_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07314__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__A1_N net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__inv_2
XANTENNA__06668__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07404_ _01719_ _01733_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nor2_1
XANTENNA__07331__B _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ net305 net335 _02562_ _03467_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07335_ top.DUT.register\[28\]\[6\] net740 net603 top.DUT.register\[5\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1061_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07266_ top.DUT.register\[29\]\[3\] net786 net595 top.DUT.register\[8\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07093__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06515__X _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ net1319 net889 _02586_ net622 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__a22o_1
X_06217_ net907 _01423_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__nor2_1
X_07197_ top.DUT.register\[10\]\[10\] net726 net756 top.DUT.register\[3\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
XANTENNA__06840__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08162__B _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout205_X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07059__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_203_Right_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_A _01534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 _04987_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_4
Xfanout521 _04981_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout532 _04963_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_4
X_09907_ _03954_ net457 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
Xfanout543 _01692_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_8
Xfanout565 net567 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_8
X_09838_ _04460_ net360 net328 top.a1.dataIn\[18\] net363 vssd1 vssd1 vccd1 vccd1
+ _04834_ sky130_fd_sc_hd__a221o_1
Xfanout587 _01564_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07553__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ top.a1.dataIn\[9\] _04766_ _04769_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_198_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11800_ _05658_ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_202_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12780_ clknet_leaf_3_clk _00326_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07305__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__A _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _05549_ _05580_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10359__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06409__Y _01526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ _05477_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ clknet_leaf_57_clk _00947_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10613_ net161 net1622 net424 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
X_11593_ _05422_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ net172 net1802 net426 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__mux2_1
X_13332_ clknet_leaf_103_clk _00878_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10094__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06831__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net186 net1488 net506 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__mux2_1
X_13263_ clknet_leaf_24_clk _00809_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ net1393 net866 net831 _06042_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13194_ clknet_leaf_118_clk _00740_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _06002_ _06005_ _06001_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10822__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07792__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _05907_ _05936_ _05921_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a21bo_1
X_11027_ net1161 _05040_ net480 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XANTENNA__09533__A1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ clknet_leaf_106_clk _00524_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09836__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ _05757_ net126 _05789_ net125 vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__o211a_1
XANTENNA__10269__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08247__B _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ top.DUT.register\[13\]\[14\] net789 _02234_ _02236_ vssd1 vssd1 vccd1 vccd1
+ _02237_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07075__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07051_ top.DUT.register\[18\]\[17\] net755 net752 top.DUT.register\[17\]\[17\] _02167_
+ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_136_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09003__A1_N _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10732__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ top.DUT.register\[24\]\[20\] net545 net627 top.DUT.register\[29\]\[20\] _03069_
+ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06904_ top.DUT.register\[13\]\[24\] net790 net774 top.DUT.register\[2\]\[24\] _02020_
+ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_182_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07884_ _02994_ _02996_ _02998_ _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__or4_1
XANTENNA__07535__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ top.pc\[29\] net853 _04637_ _04648_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06889__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ top.DUT.register\[8\]\[27\] net592 net711 top.DUT.register\[25\]\[27\] _01951_
+ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a221o_1
X_06766_ top.DUT.register\[10\]\[29\] net726 net596 top.DUT.register\[6\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
X_09554_ top.pc\[26\] _04565_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__and2_1
XANTENNA__09827__A2 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08505_ _03360_ _03612_ net281 vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__mux2_1
XANTENNA__10179__S net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09485_ _04516_ _04517_ _04518_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__a21oi_1
X_06697_ top.DUT.register\[10\]\[4\] net645 net633 top.DUT.register\[27\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout534_A _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ _02837_ _03546_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ net286 _02368_ net272 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10907__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07318_ top.DUT.register\[29\]\[7\] net787 net590 top.DUT.register\[20\]\[7\] _02434_
+ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07066__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07249_ _02356_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__nor2_8
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10260_ net251 net2279 net436 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08901__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09763__A1 _02519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10642__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net255 net1416 net441 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA__07774__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09515__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout362 _04783_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_2
Xfanout373 _04997_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_4
Xfanout384 _04978_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_6
XANTENNA__07526__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 _02521_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_2
X_12901_ clknet_leaf_39_clk _00447_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ clknet_leaf_13_clk _00378_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11086__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10089__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12763_ clknet_leaf_1_clk _00309_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ _05512_ _05556_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08635__X _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ clknet_leaf_101_clk _00240_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11645_ _05497_ _05498_ _05480_ _05488_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
XFILLER_0_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11576_ _05435_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__or2_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_1
Xinput37 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_0_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13315_ clknet_leaf_35_clk _00861_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10527_ net245 net1964 net428 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13246_ clknet_leaf_37_clk _00792_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ net267 net1909 net507 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__A _03954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10552__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ clknet_leaf_59_clk _00723_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10389_ net1561 net264 net515 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__mux2_1
XANTENNA__07765__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12128_ _05984_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12059_ _05876_ _05901_ _05907_ _05909_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07517__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire335_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ net366 net326 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13501__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ top.DUT.register\[21\]\[0\] net569 net688 top.DUT.register\[15\]\[0\] _01665_
+ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__a221o_1
XANTENNA__11077__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09270_ _04311_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07296__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06482_ net914 _01484_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nand2_4
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08221_ net298 _02175_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10727__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ net356 _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07048__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07103_ top.DUT.register\[1\]\[15\] net780 net717 top.DUT.register\[9\]\[15\] _02219_
+ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08796__A2 _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ top.DUT.register\[26\]\[17\] net681 net672 top.DUT.register\[19\]\[17\] _03199_
+ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_9_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12454__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ _02134_ _02138_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__or4_1
XANTENNA__08280__X _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10462__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06559__A1 top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ net293 _03984_ _04070_ net280 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout484_A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _01592_ _03051_ net468 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07508__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ top.DUT.register\[30\]\[27\] net695 net623 top.DUT.register\[16\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout651_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09606_ top.pc\[29\] _04622_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ top.DUT.register\[3\]\[31\] net782 net768 top.DUT.register\[11\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
X_07798_ _02908_ _02910_ _02912_ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__or4_1
XFILLER_0_210_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ _04565_ _04566_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06749_ top.DUT.register\[28\]\[28\] net739 net785 top.DUT.register\[29\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10815__A0 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ net916 top.pc\[20\] _04502_ net910 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__o211a_1
XANTENNA__07287__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ _03392_ _03398_ net287 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _04435_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__or2_1
XANTENNA__08174__Y _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07039__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11430_ _05248_ _05254_ _05257_ net478 _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a41o_2
XANTENNA__11271__A_N top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11361_ top.a1.dataIn\[27\] top.a1.dataIn\[26\] top.a1.dataIn\[28\] top.a1.dataIn\[29\]
+ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10312_ net1384 net168 net524 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__mux2_1
X_13100_ clknet_leaf_3_clk _00646_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07995__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11292_ top.a1.row1\[104\] _05149_ _05156_ _05162_ _05146_ vssd1 vssd1 vccd1 vccd1
+ _05163_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_91_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10243_ net176 net1451 net383 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
X_13031_ clknet_leaf_53_clk _00577_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10372__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07747__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A1 top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
X_10174_ net1743 net172 net526 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XANTENNA__07211__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 net1120 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_2
Xfanout181 _04867_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout192 _04841_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_1
XFILLER_0_199_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09181__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ net1125 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ clknet_leaf_24_clk _00361_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ clknet_leaf_70_clk _01320_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09121__C1 _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12746_ clknet_leaf_118_clk _00292_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07278__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10547__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ clknet_leaf_46_clk _00223_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11628_ _05454_ _05483_ _05486_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__nor3_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11559_ _05417_ _05419_ _05415_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07986__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 top.DUT.register\[9\]\[0\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold618 top.DUT.register\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold629 top.DUT.register\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09727__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ clknet_leaf_113_clk _00775_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10282__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__B2 top.pc\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ _03845_ _03858_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__nand2_1
XANTENNA__09372__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _02832_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__nand2_1
XANTENNA_wire338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09360__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _02768_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__inv_2
XANTENNA__06713__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06603_ _01607_ _01717_ _01599_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a21oi_1
X_07583_ top.DUT.register\[1\]\[15\] net705 net681 top.DUT.register\[26\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ _04362_ _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__xnor2_1
X_06534_ net746 _01647_ _01649_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__and3_1
XANTENNA__07269__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06465_ top.DUT.register\[15\]\[0\] net804 net751 top.DUT.register\[19\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a22o_1
X_09253_ _02366_ _02748_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10457__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08204_ _03318_ _03319_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__nor2_1
X_09184_ _04213_ _04216_ _04234_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor3_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06396_ _01482_ _01512_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ net829 _03251_ net468 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__o21a_1
XANTENNA__09966__A1 _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07977__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _03179_ _03180_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout699_A _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07017_ top.DUT.register\[15\]\[18\] net805 net801 top.DUT.register\[31\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
XANTENNA__10192__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__B _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09981__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__X _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13494__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13488__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ net275 _02522_ _03533_ _04050_ _01746_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__o32a_1
X_07919_ top.DUT.register\[11\]\[25\] net702 net694 top.DUT.register\[3\]\[25\] _03035_
+ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a221o_1
XFILLER_0_203_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08899_ _03009_ net459 _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10930_ net2008 net212 net485 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ net2006 net223 net489 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ clknet_leaf_37_clk _00146_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08457__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ clknet_leaf_63_clk _01121_ net1105 vssd1 vssd1 vccd1 vccd1 top.a1.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08457__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ net236 net2073 net412 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06468__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ clknet_leaf_87_clk _00077_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramstore\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10367__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12462_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[25\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11413_ _05268_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__and2_1
X_12393_ net2303 net117 _00017_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
XANTENNA__07968__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11344_ net1203 net843 _05209_ net1114 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08361__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06640__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ top.a1.row2\[16\] _05136_ _05138_ top.a1.row2\[8\] _05145_ vssd1 vssd1 vccd1
+ vccd1 _05146_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13014_ clknet_leaf_105_clk _00560_ net981 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10226_ net251 top.DUT.register\[9\]\[5\] net385 vssd1 vssd1 vccd1 vccd1 _00383_
+ sky130_fd_sc_hd__mux2_1
X_10157_ net1491 net246 net527 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XANTENNA__10830__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 top.a1.dataInTemp\[0\] vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07705__A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ net255 net1591 net389 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XANTENNA__06530__A_N top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08696__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13847_ clknet_leaf_59_clk _01370_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13778_ clknet_leaf_54_clk _01303_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07440__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06459__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ clknet_leaf_58_clk _00275_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10277__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06250_ net2239 net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[8\] sky130_fd_sc_hd__and2_1
XFILLER_0_170_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07671__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06181_ top.a1.hexop\[3\] vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07959__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 top.DUT.register\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07423__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 top.DUT.register\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold426 top.DUT.register\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 top.DUT.register\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 top.DUT.register\[14\]\[31\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ top.pc\[28\] _04622_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__and2_1
Xhold459 top.DUT.register\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap178 _05517_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_1
Xfanout906 top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ net819 _04503_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nor2_1
Xfanout917 net919 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_2
Xfanout928 net960 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_2
XFILLER_0_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload17_A clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout939 net942 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
X_08822_ _03914_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or2_1
XANTENNA__10740__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 top.DUT.register\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 top.DUT.register\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 top.DUT.register\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net318 _03848_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nand2_1
Xhold1148 top.DUT.register\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 top.DUT.register\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ net349 _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__nor2_1
X_08684_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_179_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06698__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ top.DUT.register\[26\]\[8\] net681 net542 top.DUT.register\[5\]\[8\] _02751_
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1091_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07566_ top.DUT.register\[21\]\[9\] net570 net542 top.DUT.register\[5\]\[9\] _02682_
+ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_192_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _04342_ _04346_ _04347_ net821 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06517_ _01497_ _01632_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__or2_2
XANTENNA__10187__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07497_ top.a1.instruction\[31\] net855 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09236_ _04280_ _04282_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07662__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06448_ net811 _01527_ _01528_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _04203_ _04205_ _04078_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XANTENNA__10915__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06379_ top.a1.instruction\[13\] _01489_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08118_ top.DUT.register\[1\]\[16\] net703 net663 top.DUT.register\[14\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_2_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07414__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08611__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _02928_ _02955_ _03005_ _03031_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_170_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout983_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ top.DUT.register\[31\]\[23\] net668 net548 top.DUT.register\[4\]\[23\] _03165_
+ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a221o_1
Xhold960 top.DUT.register\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 top.DUT.register\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 top.DUT.register\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net6 net862 net834 net1180 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__o22a_1
Xhold993 top.DUT.register\[5\]\[22\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net140 net1838 net453 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10650__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08127__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11962_ _05822_ _05790_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_86_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ clknet_leaf_62_clk _01234_ net1109 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[63\]
+ sky130_fd_sc_hd__dfstp_1
X_10913_ net1921 net149 net406 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11893_ _05716_ _05723_ _05753_ _05713_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12557__RESET_B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13632_ clknet_leaf_92_clk net1185 net996 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
X_10844_ net1544 net158 net495 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
XANTENNA__06428__X _01545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10097__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ clknet_leaf_0_clk _01109_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10775_ net171 net1990 net370 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12514_ clknet_leaf_93_clk _00060_ net995 vssd1 vssd1 vccd1 vccd1 top.ramstore\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09739__X _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ clknet_leaf_102_clk _01040_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06861__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12445_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[8\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10825__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13653__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12376_ top.pad.button_control.r_counter\[12\] top.pad.button_control.r_counter\[11\]
+ _06150_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_130_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11327_ top.a1.row2\[35\] _05160_ _05161_ top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1
+ _05195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13345__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _05128_ net906 net900 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ net176 net1777 net439 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
XANTENNA__10560__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net907 _01425_ _01427_ _01378_ _01420_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__o221a_1
XANTENNA__06610__Y _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_66_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08118__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06993__B _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ top.DUT.register\[2\]\[5\] net686 _02534_ _02536_ vssd1 vssd1 vccd1 vccd1
+ _02537_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07351_ _02458_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_174_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06302_ net1382 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[28\] sky130_fd_sc_hd__and2_1
XFILLER_0_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ top.DUT.register\[25\]\[2\] net712 net749 top.DUT.register\[1\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a22o_1
XANTENNA__07644__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06233_ wb.curr_state\[1\] wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__nor2_8
X_09021_ _03227_ net621 net2347 net889 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06852__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06164_ net907 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold201 top.ramaddr\[1\] vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 top.ramaddr\[24\] vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06604__B1 _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold234 top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 top.DUT.register\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 top.ramaddr\[20\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 top.DUT.register\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 top.DUT.register\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net820 _04585_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__o21ba_1
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold289 top.DUT.register\[11\]\[2\] vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 _01567_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_A _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 _01545_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_8
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_8
X_09854_ _04477_ net360 net328 top.a1.dataIn\[19\] net363 vssd1 vssd1 vccd1 vccd1
+ _04849_ sky130_fd_sc_hd__a221o_1
Xfanout747 _01645_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10470__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1104_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout769 _01560_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_2
X_08805_ _03232_ _03881_ _03261_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o21ai_1
X_09785_ top.a1.dataIn\[12\] _04766_ _04769_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_
+ sky130_fd_sc_hd__a211o_1
X_06997_ top.DUT.register\[23\]\[19\] net730 net776 top.DUT.register\[17\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout564_A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09857__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ net470 _03832_ _03833_ _02518_ _03831_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a221o_1
XFILLER_0_197_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08667_ _03723_ _03767_ net316 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__Y _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ top.DUT.register\[6\]\[11\] net577 net561 top.DUT.register\[20\]\[11\] _02734_
+ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_159_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ net320 _03658_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__or2_1
XANTENNA__07883__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _02664_ _02665_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_81_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07096__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net247 net1924 net503 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06843__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09219_ top.pc\[5\] _01809_ _04258_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a21o_1
XANTENNA__10645__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10491_ net265 net2177 net380 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ net2336 net867 net832 net129 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ _05999_ _06006_ _06010_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11112_ net96 net885 net849 net1162 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a22o_1
X_12092_ _05951_ _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_9_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 top.DUT.register\[21\]\[16\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _01400_ _01401_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nor2_1
XANTENNA__09454__B _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07020__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07571__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12994_ clknet_leaf_10_clk _00540_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11945_ _05776_ _05796_ _05797_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__and3_1
XFILLER_0_203_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _05703_ _05706_ net128 _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__a31oi_1
XANTENNA__07874__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13615_ clknet_leaf_78_clk _01156_ net1086 vssd1 vssd1 vccd1 vccd1 top.ramload\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10827_ net1426 net230 net495 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07087__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ clknet_leaf_116_clk _01092_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net246 top.DUT.register\[25\]\[6\] net373 vssd1 vssd1 vccd1 vccd1 _00896_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06834__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13477_ clknet_leaf_46_clk _01023_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13526__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ net2144 net265 net499 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09379__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ clknet_leaf_78_clk top.ru.next_FetchedData\[23\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_140_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ _06141_ _06142_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__nor2_1
XANTENNA__08051__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire365_A _02263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06920_ top.DUT.register\[16\]\[23\] net723 net754 top.DUT.register\[18\]\[23\] _02036_
+ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10290__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__A0 _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09364__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09000__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07011__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ top.DUT.register\[6\]\[26\] net597 net585 top.DUT.register\[24\]\[26\] _01967_
+ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09570_ top.pc\[27\] _04590_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__nand2_1
X_06782_ net324 _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08521_ net277 _03386_ _03395_ net271 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08452_ net285 _03561_ _03560_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07403_ net469 _02518_ _02515_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ net1275 net861 net839 _03495_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout145_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07334_ top.DUT.register\[22\]\[6\] net606 net717 top.DUT.register\[9\]\[6\] _02450_
+ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07265_ top.DUT.register\[21\]\[3\] net611 net759 top.DUT.register\[2\]\[3\] _02381_
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10465__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__RESET_B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09539__B _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout312_A _01830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _02548_ net621 net1234 net890 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06216_ _01429_ _01431_ _01432_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[0\] sky130_fd_sc_hd__or3_1
XFILLER_0_104_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ top.DUT.register\[22\]\[10\] net604 net588 top.DUT.register\[20\]\[10\] _02312_
+ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07059__B _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout500 _04995_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_4
XANTENNA_fanout681_A _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_8
X_09906_ net168 net2256 net393 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__mux2_1
Xfanout522 _04981_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_4
Xfanout544 _01689_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_4
Xfanout555 _01680_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
XANTENNA__07002__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_8
Xfanout577 net579 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_8
X_09837_ net195 net1642 net391 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__mux2_1
Xfanout588 net591 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout946_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 _01549_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_4
XANTENNA__09561__Y _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ net818 _04310_ net816 top.pc\[9\] vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_197_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07362__X _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08719_ net474 _03813_ _03815_ _02522_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_202_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _04693_ _04715_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11730_ _05586_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07856__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ _05497_ _05498_ _05473_ _05479_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a211o_1
XFILLER_0_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08905__Y _03995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13400_ clknet_leaf_38_clk _00946_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net164 net2343 net425 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07069__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11592_ _05421_ _05451_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__xor2_2
XANTENNA__08634__A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ clknet_leaf_110_clk _00877_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06816__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10375__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10543_ net174 net2089 net427 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13262_ clknet_leaf_95_clk _00808_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10474_ net188 net1731 net506 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12213_ _06048_ _05094_ net866 net1871 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13193_ clknet_leaf_27_clk _00739_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ _05994_ _05993_ _05987_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__and3b_1
XFILLER_0_20_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12075_ _05909_ _05918_ _05924_ _05908_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__or4bb_1
XANTENNA_input30_X net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net864 _05038_ _05039_ net869 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1
+ _05040_ sky130_fd_sc_hd__a32o_1
XANTENNA__07544__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13841__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07713__A _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12977_ clknet_leaf_8_clk _00523_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11928_ _05754_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nand2_1
XANTENNA__07847__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ _05683_ _05718_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_171_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06807__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13529_ clknet_leaf_58_clk _01075_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10285__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07050_ top.DUT.register\[26\]\[17\] net720 _02157_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07480__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08831__X _03924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07232__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__Y _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ top.DUT.register\[18\]\[20\] net660 net648 top.DUT.register\[12\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a22o_1
X_06903_ top.DUT.register\[18\]\[24\] net778 net777 top.DUT.register\[17\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_182_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ top.DUT.register\[26\]\[27\] net679 net552 top.DUT.register\[22\]\[27\] _02999_
+ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09622_ _01632_ _04646_ _04647_ net873 _04641_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a311o_1
X_06834_ top.DUT.register\[7\]\[27\] net707 net750 top.DUT.register\[19\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_158_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09553_ _04568_ _04574_ _04582_ _04084_ top.pc\[25\] vssd1 vssd1 vccd1 vccd1 _00106_
+ sky130_fd_sc_hd__o32a_1
X_06765_ top.DUT.register\[13\]\[29\] net788 net770 top.DUT.register\[27\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a22o_1
XANTENNA__09288__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08504_ _03507_ _03611_ net290 vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__mux2_1
XANTENNA__07299__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09484_ net916 top.pc\[21\] net911 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_210_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ top.DUT.register\[24\]\[4\] net547 net650 top.DUT.register\[12\]\[4\] _01812_
+ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ _03489_ _03545_ _02839_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ net289 _02510_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06526__X _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07317_ top.DUT.register\[11\]\[7\] net768 net709 top.DUT.register\[7\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a22o_1
XANTENNA__10195__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ net285 _03410_ _02553_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_13__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07248_ _02358_ _02360_ _02362_ _02364_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_30_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10923__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ top.DUT.register\[10\]\[11\] net726 net804 top.DUT.register\[15\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a22o_1
X_10190_ net267 net1853 net441 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06577__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
Xfanout374 _04993_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_8
Xfanout385 _04978_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
X_12900_ clknet_leaf_29_clk _00446_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_107_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ clknet_leaf_32_clk _00377_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12762_ clknet_leaf_16_clk _00308_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07829__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _05511_ _05572_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_120_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12693_ clknet_leaf_82_clk _00239_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07679__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12035__B1 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11644_ _05497_ _05498_ _05480_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a21o_1
XFILLER_0_204_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06436__X _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_1
X_11575_ top.a1.dataIn\[14\] _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and3_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XFILLER_0_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ clknet_leaf_10_clk _00860_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09747__X _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10526_ net252 net1889 net428 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__mux2_1
XANTENNA__07462__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13245_ clknet_leaf_120_clk _00791_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08006__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ net259 net1957 net507 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__mux2_1
XANTENNA__09203__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10833__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11010__A1 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07214__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ clknet_leaf_32_clk _00722_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10388_ net1475 net242 net514 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__mux2_1
XANTENNA__06568__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _05974_ _05983_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12058_ _05915_ _05916_ _05917_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ top.a1.halfData\[3\] net796 _05026_ net865 vssd1 vssd1 vccd1 vccd1 _05027_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07443__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06550_ net746 _01656_ _01662_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_47_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10824__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06481_ top.a1.instruction\[2\] _01514_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__or3b_1
XFILLER_0_28_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08151_ _01728_ _01735_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07102_ top.DUT.register\[18\]\[15\] net778 net724 top.DUT.register\[16\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XANTENNA__07453__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ top.DUT.register\[13\]\[17\] net676 net637 top.DUT.register\[25\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ _02144_ _02146_ _02147_ _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__or4_1
XANTENNA__10743__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11001__A1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06559__A2 top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ net284 _04027_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09833__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ net828 _03051_ _02618_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_149_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout477_A _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__inv_2
X_09605_ top.pc\[29\] _04622_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_162_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06817_ top.DUT.register\[20\]\[31\] net590 _01931_ _01933_ vssd1 vssd1 vccd1 vccd1
+ _01934_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07797_ top.DUT.register\[12\]\[29\] net647 net631 top.DUT.register\[27\]\[29\] _02913_
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout644_A _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06731__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ top.pc\[24\] _04534_ top.pc\[25\] vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06748_ top.DUT.register\[14\]\[28\] net794 net764 top.DUT.register\[19\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ net132 _04487_ _04501_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_210_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06679_ _01789_ _01791_ _01793_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__or4_1
XANTENNA__10918__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08484__A2 _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08418_ net277 _03527_ _03528_ net270 _03526_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__a32o_1
XANTENNA__08184__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ top.pc\[17\] _04431_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__nor2_1
X_08349_ net309 _03462_ _03433_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11360_ top.a1.dataIn\[23\] _05219_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08471__X _03581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06798__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ net2233 net170 net521 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__mux2_1
XANTENNA__10653__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ top.a1.row2\[32\] _05160_ _05161_ top.a1.row1\[112\] _05159_ vssd1 vssd1
+ vccd1 vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13030_ clknet_leaf_47_clk _00576_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10242_ net182 net1712 net384 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
X_10173_ net1632 net175 net525 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1114 net1116 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input38_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _04913_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_2
Xfanout171 _04886_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06970__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 _04867_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13863_ net1124 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11059__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ clknet_leaf_95_clk _00360_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_13794_ clknet_leaf_69_clk _01319_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12745_ clknet_leaf_26_clk _00291_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10828__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12676_ clknet_leaf_30_clk _00222_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09477__X _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _05368_ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__and2_1
XANTENNA__06789__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07986__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 top.DUT.register\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10509_ net180 net1946 net379 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
Xhold619 top.DUT.register\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10563__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11489_ _05348_ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07438__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ clknet_leaf_115_clk _00774_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13159_ clknet_leaf_56_clk _00705_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06961__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _02834_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or2_4
XANTENNA__09372__B _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _02748_ _02767_ net825 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_2
XANTENNA__06713__A2 _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ _01599_ _01718_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nand2b_4
X_07582_ top.DUT.register\[4\]\[15\] net550 net657 top.DUT.register\[28\]\[15\] _02698_
+ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09321_ _04347_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__and2_1
X_06533_ top.a1.instruction\[23\] _01648_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__or2_2
XANTENNA__10738__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09252_ _04297_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07674__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06464_ net812 _01535_ net808 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ net300 _02366_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__and2_1
X_09183_ _04213_ _04216_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06395_ net914 net913 top.a1.instruction\[6\] vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_190_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07426__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ _03241_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__nor2_2
XFILLER_0_114_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09966__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10473__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ _02047_ _03178_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07016_ net326 _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout594_A _01551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10733__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _02905_ net460 _04051_ net470 _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ top.DUT.register\[18\]\[25\] net662 net646 top.DUT.register\[10\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a22o_1
X_08898_ net398 _03005_ _03006_ net475 _03928_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_197_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ top.DUT.register\[24\]\[26\] net545 net628 top.DUT.register\[29\]\[26\] _02965_
+ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06704__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ net1865 net230 net491 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07811__A _01898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ _04538_ _04539_ _04537_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_38_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10791_ net245 net1457 net412 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__mux2_1
XANTENNA__10648__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ clknet_leaf_58_clk _00076_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramstore\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07665__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[24\] net1080 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[24\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11412_ top.a1.dataIn\[18\] _05269_ _05270_ _05271_ vssd1 vssd1 vccd1 vccd1 _05273_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07417__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net1693 net920 net38 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ top.a1.row1\[109\] _05183_ _05192_ _05206_ _05208_ vssd1 vssd1 vccd1 vccd1
+ _05209_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10383__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08361__B _03473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__A2 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ top.a1.row1\[56\] _05140_ _05142_ _05144_ net845 vssd1 vssd1 vccd1 vccd1
+ _05145_ sky130_fd_sc_hd__a2111o_1
X_13013_ clknet_leaf_101_clk _00559_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net254 net1894 net384 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XANTENNA__07196__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net1679 net252 net527 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XANTENNA__06943__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10087_ net266 net2038 net389 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
XANTENNA__08089__A _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__X _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload3_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13846_ clknet_leaf_59_clk net1152 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08160__A4 _03276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08817__A _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13777_ clknet_leaf_54_clk _01302_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _04675_ _05008_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12728_ clknet_leaf_36_clk _00274_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07120__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12659_ clknet_leaf_108_clk _00205_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06180_ wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10293__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08081__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 top.DUT.register\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__A2 _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold416 top.DUT.register\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 top.DUT.register\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold438 top.DUT.register\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06631__A1 top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold449 top.DUT.register\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout907 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_2
XFILLER_0_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _04859_ _04860_ _04861_ net816 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__o31a_1
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08384__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout929 net931 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03183_ _03913_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__nor2_1
Xhold1105 top.DUT.register\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 top.DUT.register\[21\]\[14\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 top.DUT.register\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _03848_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__inv_2
Xhold1138 top.DUT.register\[14\]\[24\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 top.DUT.register\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ net829 _02819_ net468 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08683_ _03760_ _03256_ _03252_ _02195_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09884__A1 _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ top.DUT.register\[27\]\[8\] net633 net629 top.DUT.register\[29\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
XANTENNA__07895__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10468__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ top.DUT.register\[18\]\[9\] net661 net637 top.DUT.register\[25\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09636__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09304_ _04346_ _04347_ _04342_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1084_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06516_ top.a1.instruction\[2\] _01513_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nand2_1
XANTENNA__07647__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07496_ top.a1.instruction\[31\] net855 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__nor2_2
XANTENNA__07111__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12856__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ _04280_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06447_ net809 _01550_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09166_ _04200_ _04201_ _04169_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__mux2_1
X_06378_ top.a1.instruction\[4\] net913 _01485_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__or3_2
XFILLER_0_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ top.DUT.register\[11\]\[16\] net699 net556 top.DUT.register\[8\]\[16\] _03233_
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ _01737_ _02831_ _02834_ _02847_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__and4_1
XANTENNA__08181__B _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09992__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__X _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07078__A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ top.DUT.register\[14\]\[23\] net663 net623 top.DUT.register\[16\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold950 top.DUT.register\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold961 top.DUT.register\[4\]\[27\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout976_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 top.DUT.register\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 top.DUT.register\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10931__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 top.DUT.register\[25\]\[7\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08375__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ net144 net1843 net453 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__mux2_1
X_09999_ net187 net2337 net450 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ _05787_ _05793_ _05797_ _05790_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_203_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ clknet_leaf_62_clk _01233_ net1109 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_10912_ net1432 net150 net407 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_103_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07886__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _05714_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13631_ clknet_leaf_93_clk net1195 net995 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
X_10843_ net1552 net162 net495 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10378__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13562_ clknet_leaf_15_clk _01108_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07638__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ net175 net1986 net371 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07102__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12513_ clknet_leaf_110_clk _00059_ net998 vssd1 vssd1 vccd1 vccd1 top.ramstore\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13493_ clknet_leaf_100_clk _01039_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12444_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[7\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12375_ _06151_ _06152_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11326_ top.a1.row1\[123\] _05129_ _05138_ top.a1.row2\[11\] _05193_ vssd1 vssd1
+ vccd1 vccd1 _05194_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09755__X _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ top.lcd.nextState\[5\] top.lcd.nextState\[4\] _05127_ vssd1 vssd1 vccd1 vccd1
+ _05128_ sky130_fd_sc_hd__or3_2
XANTENNA__10841__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10208_ net180 net1629 net439 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
X_11188_ net865 _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nor2_2
XANTENNA__06620__A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ net179 net1982 net443 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13829_ clknet_leaf_59_clk net1141 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.debounce_dly
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10288__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _02460_ _02462_ _02464_ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__or4_4
XFILLER_0_175_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06301_ net1285 net896 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[27\] sky130_fd_sc_hd__and2_1
XFILLER_0_127_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07281_ top.DUT.register\[5\]\[2\] net601 net751 top.DUT.register\[19\]\[2\] _02397_
+ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a221o_1
XANTENNA__08841__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09020_ net1280 net889 _03126_ net622 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__a22o_1
X_06232_ net34 net890 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_130_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06163_ net2041 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08054__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold202 top.ramstore\[28\] vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 top.DUT.register\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top.DUT.register\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06604__A1 _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 top.DUT.register\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold246 top.DUT.register\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 top.DUT.register\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 top.DUT.register\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09922_ _04590_ net361 net329 top.a1.dataIn\[26\] net364 vssd1 vssd1 vccd1 vccd1
+ _04910_ sky130_fd_sc_hd__a221o_1
Xhold279 top.DUT.register\[14\]\[8\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout704 net706 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 _01559_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_8
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_4
Xfanout737 _01531_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
XANTENNA__07626__A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ net819 _04469_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nor2_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout292_A _01774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 _01569_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_8
X_08804_ net1281 net858 net837 _03898_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__a22o_1
X_09784_ net820 _04352_ _04782_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a2bb2o_1
X_06996_ top.DUT.register\[15\]\[19\] net805 net801 top.DUT.register\[31\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XANTENNA__07580__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ net309 _03440_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__and2_1
XFILLER_0_197_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout557_A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ net322 net351 _02224_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07617_ top.DUT.register\[23\]\[11\] net565 net624 top.DUT.register\[16\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XANTENNA__10198__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ _03299_ _03304_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09987__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ net365 _02661_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07479_ top.DUT.register\[6\]\[7\] net578 net555 top.DUT.register\[22\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10926__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09218_ net918 top.pc\[5\] _04267_ top.testpc.en_latched vssd1 vssd1 vccd1 vccd1
+ _00086_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10490_ net257 net1650 net379 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08045__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _01628_ _04178_ _01598_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__o21a_1
X_12160_ _06013_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_112_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ net1225 net878 net846 top.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 _01190_
+ sky130_fd_sc_hd__a22o_1
X_12091_ _05928_ _05943_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__xor2_2
XANTENNA__10661__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold780 top.DUT.register\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 top.DUT.register\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06711__Y _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net1208 _05051_ net480 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
XANTENNA__06440__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08899__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07571__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12993_ clknet_leaf_44_clk _00539_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11104__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__B _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ _05804_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07323__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ _05703_ _05705_ net127 _05704_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_123_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10826_ net1847 net232 net495 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
X_13614_ clknet_leaf_74_clk _01155_ net1088 vssd1 vssd1 vccd1 vccd1 top.ramload\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10757_ net250 net1984 net373 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XANTENNA__10836__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13545_ clknet_leaf_28_clk _01091_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ clknet_leaf_28_clk _01022_ net1025 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10688_ net1427 net259 net498 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
X_12427_ clknet_leaf_78_clk top.ru.next_FetchedData\[22\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12358_ top.pad.button_control.r_counter\[5\] _06139_ net814 vssd1 vssd1 vccd1 vccd1
+ _06142_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10394__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ top.a1.row2\[42\] _05157_ _05174_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1
+ _05178_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10571__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ top.lcd.cnt_20ms\[13\] top.lcd.cnt_20ms\[12\] _06096_ vssd1 vssd1 vccd1 vccd1
+ _06100_ sky130_fd_sc_hd__and3_1
XANTENNA_wire358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06850_ top.DUT.register\[13\]\[26\] net789 net765 top.DUT.register\[19\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07562__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ net357 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06770__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ net462 _03626_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XANTENNA__07314__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08451_ _03318_ _03322_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__or2_1
XANTENNA__08511__B2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _01718_ _01732_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__nand2_4
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08382_ net905 top.pc\[4\] net539 _03494_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a22o_1
XANTENNA__08564__X _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07333_ top.DUT.register\[12\]\[6\] net737 net778 top.DUT.register\[18\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10746__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout138_A _04208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ top.DUT.register\[24\]\[3\] net587 net582 top.DUT.register\[4\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09003_ _01828_ net621 net1299 net891 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__a2bb2o_1
X_06215_ top.a1.hexop\[2\] top.a1.hexop\[3\] top.a1.hexop\[4\] _01428_ vssd1 vssd1
+ vccd1 vccd1 _01432_ sky130_fd_sc_hd__o31a_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08027__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ top.DUT.register\[11\]\[10\] net766 net760 top.DUT.register\[30\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06244__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A3 _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06589__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10481__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ net535 _04887_ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__and3_4
Xfanout512 _04987_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_4
Xfanout523 _04981_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout534 _04739_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_4
Xfanout545 _01689_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_4
Xfanout556 net557 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_4
X_09836_ _03800_ net455 net534 _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o211a_2
Xfanout567 _01669_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_4
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_8
Xfanout589 net591 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_4
XANTENNA__07553__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ top.DUT.register\[28\]\[20\] net738 net584 top.DUT.register\[24\]\[20\] _02095_
+ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net232 net2330 net392 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout841_A _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08718_ _01831_ _02517_ _03423_ _03371_ _03107_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__o32a_1
X_09698_ _04697_ _04700_ _04714_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08187__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07305__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__RESET_B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08649_ _03660_ _03750_ net295 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11660_ _05497_ _05498_ _05473_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ net167 net2097 net424 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10656__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_115_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11591_ _05421_ _05451_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13330_ clknet_leaf_105_clk _00876_ net982 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ net179 top.DUT.register\[18\]\[21\] net427 vssd1 vssd1 vccd1 vccd1 _00687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06435__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ clknet_leaf_113_clk _00807_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08018__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ net194 net2074 net506 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12212_ net1259 net867 net831 _06055_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__a22o_1
XANTENNA__09766__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ clknet_leaf_26_clk _00738_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ _05988_ _05995_ _05987_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10391__S net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12172__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07792__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _05908_ _05924_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__nand2_1
X_11025_ top.a1.dataInTemp\[7\] net798 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or2_1
XANTENNA__08741__B2 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06752__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__Y _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07713__B _02611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ clknet_leaf_115_clk _00522_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11927_ _05745_ _05746_ _05756_ net126 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12541__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11858_ _05683_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ net169 net1465 net413 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_106_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10566__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11789_ _05620_ _05629_ net130 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06616__Y _01733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13528_ clknet_leaf_32_clk _01074_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ clknet_leaf_108_clk _01005_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07951_ top.DUT.register\[6\]\[20\] net577 _03065_ _03067_ vssd1 vssd1 vccd1 vccd1
+ _03068_ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06902_ top.DUT.register\[14\]\[24\] net795 net590 top.DUT.register\[20\]\[24\] _02018_
+ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07882_ top.DUT.register\[2\]\[27\] net683 net635 top.DUT.register\[25\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07535__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08732__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ top.DUT.register\[22\]\[27\] net604 net784 top.DUT.register\[29\]\[27\] _01949_
+ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a221o_1
X_09621_ _04623_ _04627_ _04645_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06743__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ _01632_ _04580_ _04581_ net873 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a31o_1
X_06764_ top.DUT.register\[5\]\[29\] net600 net730 top.DUT.register\[23\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08503_ _03561_ _03610_ net315 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09483_ net132 _04503_ net916 vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06695_ top.DUT.register\[11\]\[4\] net702 net653 top.DUT.register\[17\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08434_ _02560_ _02840_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ net290 _02198_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10476__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07316_ top.DUT.register\[22\]\[7\] net606 net725 top.DUT.register\[16\]\[7\] _02432_
+ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13488__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07247_ top.DUT.register\[21\]\[8\] net610 net602 top.DUT.register\[5\]\[8\] _02363_
+ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ top.DUT.register\[16\]\[11\] net723 net593 top.DUT.register\[8\]\[11\] _02294_
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout889_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07774__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 _01799_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_167_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout364 _04768_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_2
Xfanout375 _04993_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_4
XANTENNA__07526__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
Xfanout397 _01742_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_2
X_09819_ _04808_ _04811_ _04815_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06734__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12830_ clknet_leaf_38_clk _00376_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11086__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ clknet_leaf_58_clk _00307_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _05511_ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12692_ clknet_leaf_97_clk _00238_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11643_ top.a1.dataIn\[11\] _05500_ _05502_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10386__S net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11574_ _05432_ _05433_ top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06165__A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
X_13313_ clknet_leaf_42_clk _00859_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10525_ net255 net1548 net429 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__mux2_1
X_13244_ clknet_leaf_101_clk _00790_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09739__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ net261 net1704 net507 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13175_ clknet_leaf_107_clk _00721_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08411__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _04181_ net615 _04958_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__and3_1
XANTENNA__07765__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _05952_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__xor2_1
XANTENNA__09763__X _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__inv_2
XFILLER_0_205_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07517__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ top.a1.dataInTemp\[3\] net798 vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06725__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__Y _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12959_ clknet_leaf_23_clk _00505_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06480_ top.a1.instruction\[13\] top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ _01597_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07150__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10296__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08150_ _02906_ _02931_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07101_ top.DUT.register\[22\]\[15\] net606 net762 top.DUT.register\[30\]\[15\] _02217_
+ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_151_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08081_ top.DUT.register\[3\]\[17\] net692 net668 top.DUT.register\[31\]\[17\] _03197_
+ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07032_ top.DUT.register\[8\]\[18\] net592 net580 top.DUT.register\[4\]\[18\] _02148_
+ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06803__A _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06559__A3 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ net325 net284 _01919_ _03459_ net293 vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o311a_1
XANTENNA__06964__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ _03041_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_149_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07508__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _02980_ _02981_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ top.pc\[28\] net853 _04617_ _04630_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__o22a_1
X_06816_ top.DUT.register\[16\]\[31\] net724 net772 top.DUT.register\[27\]\[31\] _01932_
+ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ top.DUT.register\[7\]\[29\] net572 net663 top.DUT.register\[14\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09535_ top.pc\[24\] top.pc\[25\] _04534_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__and3_1
X_06747_ top.DUT.register\[21\]\[28\] net609 net768 top.DUT.register\[11\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout637_A _01701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ net136 _04492_ _04500_ net823 net916 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_195_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06678_ top.DUT.register\[15\]\[1\] net689 net645 top.DUT.register\[10\]\[1\] _01794_
+ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_195_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ net290 _03385_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or2_1
X_09397_ top.pc\[17\] _04431_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout804_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__B _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ net283 _03461_ _03437_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08279_ _02111_ _02155_ net317 vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XANTENNA__10934__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13831__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ net1339 net174 net522 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__mux2_1
XANTENNA__07995__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ _05128_ _05147_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ net185 net2179 net383 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08944__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ net1781 net182 net526 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
Xfanout1104 net1111 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06955__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 net1116 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout150 net153 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 _04913_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_1
Xfanout172 _04886_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_2
Xfanout183 _04858_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
Xfanout194 _04841_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ net1123 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_199_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07380__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12813_ clknet_leaf_114_clk _00359_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13793_ clknet_leaf_70_clk _01318_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10267__A0 _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09121__A1 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12744_ clknet_leaf_25_clk _00290_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_177_Left_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07132__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12675_ clknet_leaf_33_clk _00221_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12929__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _05483_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10844__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09918__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ _05334_ _05367_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08381__Y _03494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07986__A2 _03102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold609 top.pad.button_control.r_counter\[9\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ net183 top.DUT.register\[17\]\[20\] net378 vssd1 vssd1 vccd1 vccd1 _00654_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08314__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ _05311_ _05343_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ clknet_leaf_12_clk _00773_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10439_ net1633 net196 net509 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_186_Left_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07199__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ clknet_leaf_21_clk _00704_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06946__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ top.a1.dataIn\[3\] _05965_ _05967_ _05968_ vssd1 vssd1 vccd1 vccd1 _05970_
+ sky130_fd_sc_hd__a2bb2o_1
X_13089_ clknet_leaf_43_clk _00635_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09360__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__B2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _02757_ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_195_Right_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06601_ _01602_ _01716_ _01387_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a21oi_4
X_07581_ top.DUT.register\[3\]\[15\] net693 net641 top.DUT.register\[9\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09320_ _04342_ _04346_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06532_ top.a1.instruction\[23\] _01648_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nor2_2
XFILLER_0_125_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07123__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ top.pc\[8\] _04277_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_177_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06463_ top.DUT.register\[5\]\[0\] net600 net752 top.DUT.register\[17\]\[0\] _01579_
+ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08871__B1 _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08202_ net322 _02448_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06517__B _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09182_ _04232_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06394_ _01436_ _01437_ net890 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__or3_4
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08133_ _03243_ _03245_ _03247_ _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_190_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09828__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10754__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout218_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__07977__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _02047_ _03178_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nand2_1
X_07015_ _02131_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_4__f_clk_X clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ _03928_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2_1
X_07917_ top.DUT.register\[7\]\[25\] net575 net670 top.DUT.register\[31\]\[25\] _03033_
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a221o_1
X_08897_ net270 _03826_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout754_A _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_95_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_197_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ top.DUT.register\[18\]\[26\] net660 net632 top.DUT.register\[27\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07651__X _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10929__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ top.DUT.register\[22\]\[30\] net554 net673 top.DUT.register\[19\]\[30\] _02895_
+ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07811__B _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ net133 _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nor2_1
X_10790_ net250 net1937 net413 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__mux2_1
XANTENNA__07114__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06468__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09449_ top.pc\[20\] _04467_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ clknet_leaf_78_clk top.ru.next_FetchedInstr\[23\] net1085 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[23\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _05270_ _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__and2_1
X_12391_ net1646 net920 net37 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__a21o_1
XANTENNA__10664__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06714__Y _01831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ _05188_ _05207_ _05187_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or3b_1
XANTENNA__07968__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06443__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11273_ net906 net900 top.lcd.nextState\[0\] _05143_ vssd1 vssd1 vccd1 vccd1 _05144_
+ sky130_fd_sc_hd__nor4_1
XANTENNA__06640__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10224_ net265 net1720 net384 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
X_13012_ clknet_leaf_98_clk _00558_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10155_ net2293 net253 net527 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 top.a1.dataInTemp\[5\] vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ net257 net1827 net387 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_86_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09342__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08657__X _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13845_ clknet_leaf_59_clk _01368_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10839__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_clk_X clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ clknet_leaf_64_clk _01301_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10988_ _04675_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06618__A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ clknet_leaf_107_clk _00273_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13173__RESET_B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12658_ clknet_leaf_108_clk _00204_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11609_ top.a1.dataIn\[12\] _05466_ _05467_ _05468_ vssd1 vssd1 vccd1 vccd1 _05470_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10574__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ clknet_leaf_114_clk _00135_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07959__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_194_Left_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold406 top.DUT.register\[8\]\[17\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold417 top.DUT.register\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 top.DUT.register\[18\]\[8\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 top.DUT.register\[15\]\[12\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09030__B1 _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06919__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 top.i_ready vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_55_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03183_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_14__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07592__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 top.DUT.register\[13\]\[6\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 top.DUT.register\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _02110_ _02133_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nor2_1
Xhold1128 top.DUT.register\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1139 top.DUT.register\[20\]\[29\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_77_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07702_ _02809_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08682_ net1336 net858 net837 _03782_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a22o_1
XANTENNA__07344__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_179_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07633_ top.DUT.register\[3\]\[8\] net693 net550 top.DUT.register\[4\]\[8\] _02749_
+ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a221o_1
XANTENNA__06698__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ top.DUT.register\[20\]\[9\] net562 net546 top.DUT.register\[24\]\[9\] _02680_
+ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06528__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ net347 _04345_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__or2_1
X_06515_ top.a1.instruction\[2\] _01482_ _01512_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__and3_4
XFILLER_0_76_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07495_ _02438_ _02447_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__or3_4
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1077_A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ top.pc\[6\] _02528_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a21o_1
X_06446_ net809 _01562_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ net822 _04216_ _04217_ _04171_ net400 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__o32a_1
XANTENNA__06870__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10484__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__B _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06377_ net913 _01485_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout502_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08116_ top.DUT.register\[20\]\[16\] net560 net647 top.DUT.register\[12\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a22o_1
X_09096_ _02561_ _02797_ _02844_ _03104_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08047_ top.DUT.register\[6\]\[23\] net576 net699 top.DUT.register\[11\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold940 top.DUT.register\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 top.DUT.register\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09001__A1_N _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold962 top.DUT.register\[10\]\[18\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 top.DUT.register\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06550__X _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold984 top.DUT.register\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 top.DUT.register\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__B _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net191 net2003 net450 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07583__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _02932_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09016__A1_N _03202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08127__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _05783_ _05806_ _05814_ _05819_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__or4b_1
XANTENNA__07335__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ net1583 net157 net406 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__mux2_1
XANTENNA__07886__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _05708_ net128 _05707_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ clknet_leaf_92_clk net1199 net996 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
X_10842_ net1862 net166 net496 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13561_ clknet_leaf_56_clk _01107_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10773_ net182 net2099 net372 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12512_ clknet_leaf_75_clk _00058_ net1084 vssd1 vssd1 vccd1 vccd1 top.ramstore\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13492_ clknet_leaf_103_clk _01038_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[6\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[6\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_23_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10394__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06861__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12374_ net1433 _06150_ net814 vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ top.a1.row2\[3\] _05132_ _05136_ top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1
+ _05193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ top.lcd.nextState\[1\] top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05127_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ net186 net2031 net439 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
X_11187_ _05012_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nand2_1
XANTENNA__06620__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A1_N net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ net184 net1478 net443 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12411__Q top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ net190 net1601 net446 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09866__A2 _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10569__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06619__Y _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13828_ clknet_leaf_59_clk _00017_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.noisy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13759_ clknet_leaf_65_clk _01284_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08834__Y _03927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06300_ net2346 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[26\] sky130_fd_sc_hd__and2_1
X_07280_ top.DUT.register\[14\]\[2\] net793 net585 top.DUT.register\[24\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06231_ top.ru.state\[6\] top.busy_o top.ru.state\[3\] vssd1 vssd1 vccd1 vccd1 _01438_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06852__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06162_ top.lcd.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__09946__X _04932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 top.DUT.register\[31\]\[5\] vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 top.DUT.register\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06604__A2 _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 top.ramaddr\[31\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold236 top.DUT.register\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold247 top.DUT.register\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 top.DUT.register\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 top.DUT.register\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _04898_ _04906_ _04907_ _04191_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 net706 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_8
Xfanout716 _01559_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_4
X_09852_ _04842_ _04845_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__xnor2_1
Xfanout727 _01544_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
Xfanout738 net741 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
XANTENNA__07565__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 _01586_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
XANTENNA__06530__B top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ net903 top.pc\[22\] net539 _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09783_ _01594_ _04784_ net362 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a21o_1
X_06995_ _02070_ _02111_ net318 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout285_A _01800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08734_ net309 _03462_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__and2_1
XANTENNA__07317__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10479__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _01729_ _03253_ _03256_ net459 _03763_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout452_A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ top.DUT.register\[14\]\[11\] net664 net545 top.DUT.register\[24\]\[11\] _02732_
+ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a221o_1
X_08596_ _03503_ _03569_ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a21o_1
XANTENNA__09609__A2 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ net365 _02661_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08293__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07096__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ top.DUT.register\[11\]\[7\] net701 net677 top.DUT.register\[13\]\[7\] _02594_
+ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09217_ net133 _04256_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06843__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06429_ net811 _01524_ net808 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09856__X _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _01628_ _04177_ _04198_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09793__A1 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10942__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _03424_ _03464_ _03505_ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11110_ net1313 net883 net848 top.ramstore\[28\] vssd1 vssd1 vccd1 vccd1 _01189_
+ sky130_fd_sc_hd__a22o_1
X_12090_ _05938_ _05944_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__xnor2_1
Xhold770 top.DUT.register\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 top.DUT.register\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ net864 _05049_ _05050_ net869 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1
+ _05051_ sky130_fd_sc_hd__a32o_1
Xhold792 top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06440__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07308__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ clknet_leaf_14_clk _00538_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07552__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11943_ _05799_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nand2_1
XANTENNA__10389__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11874_ _05732_ _05733_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_123_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ clknet_leaf_78_clk _01154_ net1087 vssd1 vssd1 vccd1 vccd1 top.ramload\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10825_ net1770 net238 net495 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09479__A _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ clknet_leaf_31_clk _01090_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10756_ net254 net1895 net373 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13475_ clknet_leaf_35_clk _01021_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06834__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ net2180 net262 net499 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XANTENNA__06615__B _01727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__X _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ clknet_leaf_78_clk top.ru.next_FetchedData\[21\] net1085 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__Q top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ top.pad.button_control.r_counter\[5\] top.pad.button_control.r_counter\[4\]
+ _06137_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__and3_1
XANTENNA__10852__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ top.a1.row2\[18\] _05136_ _05149_ top.a1.row1\[106\] _05142_ vssd1 vssd1
+ vccd1 vccd1 _05177_ sky130_fd_sc_hd__a221o_1
X_12288_ top.lcd.cnt_20ms\[12\] top.lcd.cnt_20ms\[11\] _06095_ top.lcd.cnt_20ms\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__a31o_1
X_11239_ net871 _05032_ _05044_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07011__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06780_ _01891_ _01894_ _01895_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__nor4_1
XFILLER_0_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10299__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ net315 _03506_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07401_ _01718_ _01732_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__and2_4
X_08381_ net462 _03468_ _03492_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08732__A1_N net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07332_ net297 _02448_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07263_ top.DUT.register\[14\]\[3\] net795 net713 top.DUT.register\[25\]\[3\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a221o_1
XANTENNA__06825__A2 _01941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06214_ top.a1.hexop\[3\] _01428_ _01431_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[7\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ net1263 net889 _01854_ net622 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07194_ top.DUT.register\[28\]\[10\] net738 net758 top.DUT.register\[2\]\[10\] _02310_
+ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08578__A2 _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10762__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout200_A _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07250__A2 _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ net817 _04893_ _04889_ _04888_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a211o_1
Xfanout502 net504 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_8
Xfanout513 net516 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_6
Xfanout524 _04981_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_4
XANTENNA__07538__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06260__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
Xfanout546 _01689_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07002__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _04829_ _04830_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__or3_1
Xfanout557 _01677_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_4
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 _01651_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_4
XANTENNA_fanout667_A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _03603_ net456 net535 _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o211a_2
X_06978_ top.DUT.register\[23\]\[20\] net730 net767 top.DUT.register\[11\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
XANTENNA__07372__A _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net398 _03104_ _03105_ net475 _03765_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__o221a_1
X_09697_ _04699_ _04701_ _04694_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_197_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout834_A _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08187__B _02305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09998__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ _03701_ _03749_ net320 vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__mux2_1
XANTENNA__10002__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08579_ net312 _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nand2_1
XANTENNA__10937__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10610_ net170 net2047 net422 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
XANTENNA__07069__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _05432_ _05433_ _05414_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net185 net1467 net427 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06816__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13610__Q top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06435__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13260_ clknet_leaf_116_clk _00806_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ net195 net2134 net505 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12211_ net2208 net866 net831 _06063_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__a22o_1
XANTENNA__09766__A1 _03603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10672__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ clknet_leaf_49_clk _00737_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07777__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ _05994_ _05993_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07241__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06451__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ _05932_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__and2_1
XANTENNA__07529__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__X _02951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ top.a1.data\[3\] net796 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or2_1
XANTENNA__09762__A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11089__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12975_ clknet_leaf_22_clk _00521_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11926_ _05785_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12492__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11857_ _05674_ _05677_ _05687_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__o21a_1
XANTENNA__10847__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ net171 net2147 net410 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__mux2_1
XANTENNA__08257__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ _05640_ _05646_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_171_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13527_ clknet_leaf_111_clk _01073_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06807__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ net185 net2254 net415 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07480__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ clknet_leaf_107_clk _01004_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ clknet_leaf_54_clk top.ru.next_FetchedData\[4\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10582__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__clkbuf_4
X_13389_ clknet_leaf_113_clk _00935_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07768__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07232__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09509__A1 _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ top.DUT.register\[20\]\[20\] net561 net624 top.DUT.register\[16\]\[20\] _03066_
+ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a221o_1
X_06901_ top.DUT.register\[5\]\[24\] net602 net768 top.DUT.register\[11\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
X_07881_ top.DUT.register\[6\]\[27\] net576 net631 top.DUT.register\[27\]\[27\] _02997_
+ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_182_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _04623_ _04627_ _04645_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__o21ai_2
X_06832_ top.DUT.register\[12\]\[27\] net734 net758 top.DUT.register\[2\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09551_ _04558_ _04562_ _04579_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__or3_1
X_06763_ top.DUT.register\[15\]\[29\] net804 net800 top.DUT.register\[31\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08502_ _03306_ _03319_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__or2_1
XANTENNA__09142__C1 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07299__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09482_ net136 _04508_ _04515_ net821 vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__o22a_1
X_06694_ top.DUT.register\[21\]\[4\] net570 net665 top.DUT.register\[14\]\[4\] _01810_
+ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08496__B2 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08433_ _03539_ _03540_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__and3_1
XANTENNA__10757__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08364_ net289 _02286_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nand2_1
XANTENNA__09445__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ top.DUT.register\[28\]\[7\] net740 net599 top.DUT.register\[6\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
X_08295_ _02408_ _02429_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout415_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ top.DUT.register\[11\]\[8\] net768 net590 top.DUT.register\[20\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ top.DUT.register\[14\]\[11\] net793 net581 top.DUT.register\[4\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22o_1
XANTENNA__10492__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout784_A _01534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07086__B net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_167_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 net323 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout376 _04993_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_8
X_09818_ _04808_ _04811_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__and3_1
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_6
Xfanout398 _01742_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
XANTENNA__07931__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09749_ net820 _04275_ top.a1.dataIn\[6\] net813 vssd1 vssd1 vccd1 vccd1 _04757_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_179_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ clknet_leaf_32_clk _00306_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11711_ _05512_ _05535_ _05541_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10294__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10667__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12691_ clknet_leaf_111_clk _00237_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11642_ _05500_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__and2_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_1
X_13312_ clknet_leaf_14_clk _00858_ net980 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_1
X_10524_ net267 net1839 net429 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07462__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__A1 _03465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ clknet_leaf_5_clk _00789_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ net242 net1995 net505 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ clknet_leaf_105_clk _00720_ net981 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07214__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__B2 _03522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386_ net1383 net140 net433 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__mux2_1
X_12125_ _05972_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__and2_1
XANTENNA__08962__A2 _03967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09492__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ _05869_ _05902_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ net1173 _05025_ _05013_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07922__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ clknet_leaf_37_clk _00504_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10577__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ clknet_leaf_42_clk _00435_ net1071 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11262__A top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_116_clk_X clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07100_ top.DUT.register\[3\]\[15\] net782 net768 top.DUT.register\[11\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_151_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08080_ top.DUT.register\[15\]\[17\] net688 net656 top.DUT.register\[28\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a22o_1
XANTENNA__07453__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08571__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07031_ top.DUT.register\[12\]\[18\] net734 net600 top.DUT.register\[5\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07205__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08982_ _02881_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ _03043_ _03045_ _03047_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_149_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout198_A _04833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _01981_ _02978_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and2_1
XANTENNA__06716__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09603_ net136 _04620_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__o21ai_1
X_06815_ top.DUT.register\[14\]\[31\] net794 net786 top.DUT.register\[29\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ top.DUT.register\[24\]\[29\] net544 net659 top.DUT.register\[18\]\[29\] _02911_
+ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09534_ top.pc\[24\] _04084_ _04549_ _04564_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06746_ top.DUT.register\[12\]\[28\] net735 net605 top.DUT.register\[22\]\[28\] _01862_
+ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _04497_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_195_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06677_ top.DUT.register\[9\]\[1\] net641 net626 top.DUT.register\[16\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12432__RESET_B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08416_ net286 _03387_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__or2_1
X_09396_ _01415_ net853 net873 _04434_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06266__A top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ _03438_ _03460_ net287 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08278_ net287 _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06553__X _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13638__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06652__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ _02340_ _02345_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__nor2_8
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09864__X _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ net190 net2092 net382 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12504__Q top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net1900 net184 net526 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__10950__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13220__RESET_B net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1105 net1107 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1116 net1120 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout140 net142 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_2
Xfanout151 net153 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout162 net165 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
Xfanout173 _04886_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_1
Xfanout184 _04858_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_98_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07904__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 net198 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
X_13861_ net1122 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_198_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12812_ clknet_leaf_115_clk _00358_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13792_ clknet_leaf_70_clk _01317_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ clknet_leaf_56_clk _00289_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08501__A1_N net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10397__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06176__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12674_ clknet_leaf_12_clk _00220_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06891__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ _05484_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13656__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _05395_ _05396_ _05397_ net248 vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10507_ net189 net2313 net378 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11487_ _05315_ _05335_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13226_ clknet_leaf_117_clk _00772_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09774__X _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10438_ net2051 net201 net509 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12414__Q top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13157_ clknet_leaf_47_clk _00703_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10860__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ net1835 net209 net430 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12108_ _05967_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nand2_1
X_13088_ clknet_leaf_13_clk _00634_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ _05878_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08699__A1 _02519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06600_ _01387_ _01603_ _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__or3_2
X_07580_ top.DUT.register\[6\]\[15\] net578 net661 top.DUT.register\[18\]\[15\] _02696_
+ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06531_ top.a1.instruction\[22\] net799 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10100__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ top.pc\[8\] _04277_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__and2_1
X_06462_ top.DUT.register\[14\]\[0\] net793 net720 top.DUT.register\[26\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07674__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ net285 _03313_ _03316_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a21o_1
XANTENNA__06882__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06393_ net1284 net1141 _01510_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _01834_ net344 vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08132_ top.DUT.register\[21\]\[16\] net568 net659 top.DUT.register\[18\]\[16\] _03248_
+ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07469__X _02586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07426__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08505__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07188__Y _02305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ _02048_ _03178_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__and2_2
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07014_ _02129_ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10770__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08240__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ net477 _02903_ _02904_ net398 vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout482_A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ top.DUT.register\[26\]\[25\] net681 net559 top.DUT.register\[8\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ net311 _03663_ _03985_ net280 vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_166_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07847_ top.DUT.register\[9\]\[26\] net640 _02963_ vssd1 vssd1 vccd1 vccd1 _02964_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_197_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07778_ top.DUT.register\[15\]\[30\] net689 net657 top.DUT.register\[28\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ top.pc\[24\] _04534_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06729_ top.DUT.register\[12\]\[3\] net650 net629 top.DUT.register\[29\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08195__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10010__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ net916 top.pc\[19\] _04483_ net910 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07665__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06873__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__Y _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ _01414_ net853 net873 _04418_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__o22ai_1
XANTENNA__10945__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11410_ top.a1.dataIn\[19\] _05243_ net479 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or3b_1
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12390_ net2087 net920 net36 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__a21o_1
XANTENNA__07417__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ top.a1.row1\[13\] _05127_ _05152_ _05140_ top.a1.row1\[61\] vssd1 vssd1 vccd1
+ vccd1 _05207_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06443__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11272_ top.lcd.nextState\[5\] top.lcd.nextState\[4\] top.lcd.nextState\[1\] vssd1
+ vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or3b_1
X_13011_ clknet_leaf_94_clk _00557_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ net258 net2141 net384 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XANTENNA__10680__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10154_ net1423 net265 net527 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10085_ net263 top.DUT.register\[5\]\[1\] net388 vssd1 vssd1 vccd1 vccd1 _00251_
+ sky130_fd_sc_hd__mux2_1
Xhold7 top.a1.dataInTemp\[1\] vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
X_13844_ clknet_leaf_59_clk _01367_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12229__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06458__X _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ clknet_leaf_61_clk _01300_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10987_ _00017_ _01426_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ clknet_leaf_102_clk _00272_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12409__Q top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10855__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12657_ clknet_leaf_9_clk _00203_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11608_ _05467_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__and2_1
XANTENNA__08605__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08605__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ clknet_leaf_3_clk _00134_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11539_ _05371_ _05374_ _05379_ _05399_ _05380_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__a41o_1
XANTENNA__08081__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 top.DUT.register\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 top.DUT.register\[22\]\[6\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold429 top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13209_ clknet_leaf_61_clk _00755_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10590__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout909 top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_55_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07041__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _03082_ net460 _03843_ net471 _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__a221o_1
Xhold1107 top.DUT.register\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 top.DUT.register\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 top.DUT.register\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ _02811_ _02813_ _02815_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__or4_1
X_08681_ net902 top.pc\[16\] net537 _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07632_ top.DUT.register\[14\]\[8\] net665 net641 top.DUT.register\[9\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_179_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07563_ top.DUT.register\[28\]\[9\] net657 net633 top.DUT.register\[27\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
X_09302_ net347 _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ top.a1.instruction\[7\] _01486_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_192_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07494_ _02591_ _02610_ net826 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_4
XANTENNA__07647__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ top.pc\[6\] _02528_ _04268_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__o21a_1
XANTENNA__06855__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06445_ _01520_ _01524_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ _04212_ _04215_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nor2_1
X_06376_ top.lcd.cnt_500hz\[13\] _01496_ top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1
+ vccd1 top.lcd.lcd_en sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _03229_ _03230_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__and2_2
XANTENNA__10403__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09095_ _02904_ _02981_ _03844_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__and3_1
XANTENNA__08072__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06263__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ top.DUT.register\[18\]\[23\] net659 net631 top.DUT.register\[27\]\[23\] _03162_
+ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a221o_1
XANTENNA__07280__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 top.DUT.register\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 top.DUT.register\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold952 top.DUT.register\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 top.DUT.register\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold974 top.DUT.register\[28\]\[16\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__B2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 top.DUT.register\[20\]\[8\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 top.DUT.register\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08375__A3 _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07032__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A2 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ net195 net2244 net451 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10005__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _02954_ _04013_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__nand2b_1
X_08879_ net312 _03636_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10910_ net1961 net158 net407 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__inv_2
XANTENNA__07886__A2 _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ top.DUT.register\[27\]\[23\] net170 net493 vssd1 vssd1 vccd1 vccd1 _00977_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09088__A1 _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07099__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ clknet_leaf_33_clk _01106_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10772_ net183 net1425 net371 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XANTENNA__07638__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ clknet_leaf_89_clk _00057_ net1015 vssd1 vssd1 vccd1 vccd1 top.ramstore\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06846__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ clknet_leaf_108_clk _01037_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10675__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ clknet_leaf_54_clk top.ru.next_FetchedInstr\[5\] net1077 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12373_ top.pad.button_control.r_counter\[11\] _06150_ vssd1 vssd1 vccd1 vccd1 _06151_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11324_ net845 _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__or2_1
XANTENNA__07271__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__X _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ net1296 net403 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_26_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10206_ net187 net2334 net438 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
XANTENNA__07023__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _04676_ net870 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nand2_2
X_10137_ net187 net1913 net442 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
XANTENNA__09753__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ net191 net2247 net447 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13827_ clknet_leaf_60_clk _01352_ net1102 vssd1 vssd1 vccd1 vccd1 top.pad.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_35_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09768__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ clknet_leaf_65_clk _01283_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12709_ clknet_leaf_40_clk _00255_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10585__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09659__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ clknet_leaf_79_clk _00005_ net1085 vssd1 vssd1 vccd1 vccd1 top.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06230_ net34 _01437_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06161_ top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08054__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 top.DUT.register\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 top.a1.row1\[18\] vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 top.DUT.register\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold237 top.a1.row1\[56\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 top.DUT.register\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _04898_ _04907_ _04906_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__o21a_1
Xhold259 top.DUT.register\[27\]\[2\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 _01654_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ _04845_ _04842_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nand2b_1
Xfanout717 _01559_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_8
Xfanout728 _01544_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_8
Xfanout739 net741 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
X_08802_ _02518_ _03883_ _03892_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a211o_1
X_09782_ top.pc\[12\] _04359_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ net299 _02089_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a21o_1
X_08733_ _03764_ _03829_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout180_A _04867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09711__C1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__inv_2
XANTENNA__07868__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06539__A top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ top.DUT.register\[17\]\[11\] net652 net628 top.DUT.register\[29\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11164__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ net280 _03498_ _03501_ net269 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a22o_1
XANTENNA__06258__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _02264_ _02661_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06828__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08293__A2 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ top.DUT.register\[3\]\[7\] net693 net661 top.DUT.register\[18\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ net137 _04258_ _04259_ _04265_ net918 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06428_ net812 _01524_ net808 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__and3_2
XFILLER_0_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ _01628_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06359_ top.a1.instruction\[3\] _01481_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__nor2_2
XANTENNA__08045__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ net279 _03503_ _04008_ _04129_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09793__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08029_ top.DUT.register\[19\]\[19\] net671 net635 top.DUT.register\[25\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a22o_1
Xhold760 top.DUT.register\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 top.DUT.register\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 top.DUT.register\[29\]\[29\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09872__X _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ top.a1.dataInTemp\[11\] net798 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold793 top.DUT.register\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10560__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12991_ clknet_leaf_31_clk _00537_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ _05785_ _05796_ _05797_ _05772_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a31o_1
XANTENNA__07552__B _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11873_ _05732_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ clknet_leaf_74_clk _01153_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramload\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10824_ net2165 net245 net495 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13543_ clknet_leaf_53_clk _01089_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06819__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ net267 net1639 net372 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09479__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13474_ clknet_leaf_11_clk _01020_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08951__X _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ net1908 net241 net498 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_80_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09769__C1 _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12425_ clknet_leaf_78_clk top.ru.next_FetchedData\[20\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07244__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _06139_ _06140_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11307_ top.a1.row1\[58\] _05140_ _05158_ top.a1.row1\[10\] _05175_ vssd1 vssd1 vccd1
+ vccd1 _05176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12287_ net1190 _06096_ _06098_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11238_ _05119_ net1266 net402 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12422__Q top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ net924 net1283 net877 _05084_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11265__A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06770__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07400_ _01735_ _01744_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__or2_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ _03474_ _03481_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ _02438_ _02447_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__nor2_4
XFILLER_0_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07262_ top.DUT.register\[9\]\[3\] net718 net762 top.DUT.register\[30\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09001_ _01773_ net621 net1159 net890 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__a2bb2o_1
X_06213_ top.a1.halfData\[0\] _01430_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_154_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09015__A1_N _03251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08027__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07193_ top.DUT.register\[14\]\[10\] net792 net752 top.DUT.register\[17\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07235__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06589__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _04890_ _04891_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__xnor2_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_6
Xfanout514 net516 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_4
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout536 _04739_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
Xfanout547 _01689_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
X_09834_ _04445_ net362 net329 top.a1.dataIn\[17\] net364 vssd1 vssd1 vccd1 vccd1
+ _04831_ sky130_fd_sc_hd__a221o_1
Xfanout558 _01677_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_8
Xfanout569 _01666_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_206_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__A _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ top.a1.dataIn\[8\] _04766_ _04769_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_198_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06977_ top.DUT.register\[27\]\[20\] net771 net765 top.DUT.register\[19\]\[20\] _02093_
+ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout562_A _01673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ net303 _03405_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__or2_1
XANTENNA__07372__B _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _04692_ _04698_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08647_ _03296_ _03300_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ net282 _03485_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07529_ top.DUT.register\[21\]\[13\] net568 net548 top.DUT.register\[4\]\[13\] _02645_
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ net187 top.DUT.register\[18\]\[19\] net426 vssd1 vssd1 vccd1 vccd1 _00685_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10953__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ net201 net2068 net505 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ net1373 net866 net831 _06068_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07226__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__B2 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ clknet_leaf_49_clk _00736_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09766__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ _05995_ _05999_ _05996_ _05988_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_94_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06451__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12072_ _05898_ _05926_ _05929_ _05881_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__or4b_1
Xhold590 top.DUT.register\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net1166 _05037_ _05013_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06752__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ clknet_leaf_97_clk _00520_ net1001 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06179__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ _05767_ _05768_ _05772_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11856_ _05703_ _05706_ _05708_ _05715_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a211o_1
XANTENNA__06907__A _02023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ net176 net1695 net411 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_109_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11787_ _05609_ _05642_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_171_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10738_ net187 net2160 net414 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
X_13526_ clknet_leaf_104_clk _01072_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07465__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12417__Q top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10863__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_7_clk _01003_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ net199 net2280 net418 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12408_ clknet_leaf_54_clk top.ru.next_FetchedData\[3\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07217__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_3_clk _00934_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12550__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ top.pad.count\[0\] net920 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09509__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06900_ top.DUT.register\[19\]\[24\] net764 _02014_ _02016_ vssd1 vssd1 vccd1 vccd1
+ _02017_ sky130_fd_sc_hd__a211o_1
X_07880_ top.DUT.register\[7\]\[27\] net572 net540 top.DUT.register\[5\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a22o_1
XANTENNA__08569__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13756__RESET_B net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ top.DUT.register\[21\]\[27\] net608 net752 top.DUT.register\[17\]\[27\] _01947_
+ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06743__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ _04558_ _04562_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10103__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ net324 _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__nand2_1
X_08501_ net396 _02691_ _02690_ net476 vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07760__X _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09481_ _04509_ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06693_ top.DUT.register\[13\]\[4\] net677 net642 top.DUT.register\[9\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08432_ net394 _03535_ _03542_ net469 vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__a22oi_1
XANTENNA__07920__B net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ _02518_ _03475_ _03474_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07314_ top.DUT.register\[14\]\[7\] net794 net583 top.DUT.register\[4\]\[7\] _02430_
+ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a221o_1
XANTENNA__07456__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _02845_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08591__X _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07245_ top.DUT.register\[23\]\[8\] net732 net764 top.DUT.register\[19\]\[8\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a221o_1
XANTENNA__10773__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06823__Y _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07176_ top.DUT.register\[21\]\[11\] net609 net712 top.DUT.register\[25\]\[11\] _02292_
+ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08956__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 _01711_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_167_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout777_A _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
Xfanout377 _04993_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
X_09817_ top.pc\[16\] _04425_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__xnor2_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_6
Xfanout399 _01742_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08198__B _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ net250 net1906 net392 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09679_ top.pad.keyCode\[1\] top.pad.keyCode\[2\] top.pad.keyCode\[3\] top.pad.keyCode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or4b_2
XANTENNA__10948__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _05549_ _05551_ _05553_ _05563_ _05569_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__a311o_2
X_12690_ clknet_leaf_115_clk _00236_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07695__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11641_ top.a1.dataIn\[12\] _05497_ _05498_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11572_ _05378_ _05428_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13311_ clknet_leaf_32_clk _00857_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10523_ net260 net1883 net427 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
XANTENNA__10683__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ clknet_leaf_15_clk _00788_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09739__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ net614 _04729_ _04738_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__or3_4
XFILLER_0_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13173_ clknet_leaf_81_clk _00719_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10385_ net2175 net145 net432 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12124_ _05977_ _05980_ _05970_ _05974_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a211o_1
X_12055_ _05891_ _05910_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__xnor2_1
X_11006_ top.a1.dataIn\[2\] net869 _05022_ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06725__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10858__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ clknet_leaf_119_clk _00503_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08836__B _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ _05739_ _05744_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__nor2_1
XANTENNA__07686__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ clknet_leaf_35_clk _00434_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06637__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ top.a1.dataIn\[6\] _05697_ _05698_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13509_ clknet_leaf_40_clk _01055_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10593__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07030_ top.DUT.register\[13\]\[18\] net788 net754 top.DUT.register\[18\]\[18\] _02135_
+ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_180_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _02905_ _04057_ _02903_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06964__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ top.DUT.register\[12\]\[25\] net649 net641 top.DUT.register\[9\]\[25\] _03048_
+ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_149_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08299__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__inv_2
XANTENNA__12224__A2_N _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06814_ top.DUT.register\[15\]\[31\] net806 net802 top.DUT.register\[31\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a22o_1
X_09602_ _04627_ _04628_ net873 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o21ba_1
X_07794_ top.DUT.register\[9\]\[29\] net639 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09533_ _01632_ _04563_ _04555_ net873 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a211o_1
X_06745_ top.DUT.register\[5\]\[28\] net601 net776 top.DUT.register\[17\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a22o_1
XANTENNA__10768__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A _04747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08746__B _03473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09464_ _04479_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06676_ top.DUT.register\[11\]\[1\] net701 net558 top.DUT.register\[8\]\[1\] _01792_
+ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_195_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07141__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ net290 _03394_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11172__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ net135 _04423_ _04433_ net131 _04430_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout525_A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout146_X net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07429__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08277_ net284 _02026_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07228_ _02332_ _02342_ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__or3_2
XFILLER_0_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ top.DUT.register\[29\]\[12\] net784 net707 top.DUT.register\[7\]\[12\] _02275_
+ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a221o_1
XANTENNA__10008__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10170_ net1505 net188 net525 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06955__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_2
Xfanout130 _05649_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_2
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout163 net165 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 _04878_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_2
Xfanout185 _04858_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
X_13860_ top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07380__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ clknet_leaf_6_clk _00357_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10678__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13791_ clknet_leaf_70_clk _01316_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12742_ clknet_leaf_19_clk _00288_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07132__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12673_ clknet_leaf_45_clk _00219_ net1066 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11624_ _05449_ _05465_ _05450_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_13_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08093__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ _05395_ net248 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_42_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10506_ net191 net2126 net378 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11486_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13225_ clknet_leaf_9_clk _00771_ net973 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net1492 net205 net511 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07199__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13156_ clknet_leaf_28_clk _00702_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10368_ net1796 net213 net430 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06946__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ _05898_ _05963_ _05957_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13087_ clknet_leaf_31_clk _00633_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ net1879 net221 net522 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
X_12038_ _05892_ _05894_ _05882_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09950__B _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10588__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09648__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ top.a1.instruction\[20\] top.a1.instruction\[21\] _01644_ vssd1 vssd1 vccd1
+ vccd1 _01647_ sky130_fd_sc_hd__and3b_2
XFILLER_0_29_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07123__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06461_ net811 _01518_ net808 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ net313 _03314_ _03315_ net286 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ _01834_ net344 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nor2_1
X_06392_ _01503_ _01507_ _01508_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ top.DUT.register\[31\]\[16\] net667 net651 top.DUT.register\[17\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ _02048_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07831__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07013_ _02113_ _02116_ _02118_ _02120_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13771__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06937__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ net275 _03532_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nor2_1
X_07915_ _03030_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nor2_2
X_08895_ _03907_ _03984_ net293 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07846_ top.DUT.register\[1\]\[26\] net704 net656 top.DUT.register\[28\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a22o_1
XANTENNA__07898__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07777_ top.DUT.register\[3\]\[30\] net693 net650 top.DUT.register\[12\]\[30\] _02893_
+ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a221o_1
XANTENNA__10498__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout642_A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06728_ top.DUT.register\[30\]\[3\] net697 net677 top.DUT.register\[13\]\[3\] _01844_
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a221o_1
X_09516_ _01416_ net853 net873 _04547_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08311__B2 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ net131 _04469_ _04482_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06659_ _01630_ _01638_ _01748_ net400 net856 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_42_clk_X clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09378_ net135 _04407_ _04417_ net131 _04416_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12848__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _02848_ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11340_ top.a1.row1\[101\] _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07822__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11271_ top.lcd.nextState\[1\] top.lcd.nextState\[0\] top.a1.row2\[12\] _05141_ vssd1
+ vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and4b_1
XANTENNA__10961__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13010_ clknet_leaf_106_clk _00556_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10222_ net261 net1445 net385 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XANTENNA__07836__A _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06740__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ net1458 net257 net526 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09327__B1 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net240 net2088 net386 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
Xhold8 top.a1.dataInTemp\[6\] vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06739__X _01856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09115__X _04168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__A2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ clknet_leaf_59_clk _01366_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06561__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10201__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ net920 _01421_ _01426_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or4b_1
X_13774_ clknet_leaf_67_clk _01299_ net1114 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ clknet_leaf_83_clk _00271_ net1007 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12656_ clknet_leaf_115_clk _00202_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ top.a1.dataIn\[13\] _05437_ net207 vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12587_ clknet_leaf_6_clk _00133_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11538_ _05389_ _05394_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 top.DUT.register\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold419 top.DUT.register\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10871__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11469_ _05322_ _05329_ _05320_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a21o_2
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13208_ clknet_leaf_37_clk _00754_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06919__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_111_clk _00685_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 top.DUT.register\[4\]\[18\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 top.DUT.register\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ top.DUT.register\[20\]\[12\] net560 net627 top.DUT.register\[29\]\[12\] _02816_
+ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a221o_1
XFILLER_0_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ net463 _03761_ _03774_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a211o_1
XANTENNA__08577__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07344__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__B2 _03647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ top.a1.instruction\[29\] _01613_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_205_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10111__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ top.DUT.register\[15\]\[9\] net690 net669 top.DUT.register\[31\]\[9\] _02678_
+ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a221o_1
X_09301_ net854 _01635_ net619 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06513_ net841 net401 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_192_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07493_ _02600_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ top.pc\[7\] _02566_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__xnor2_1
X_06444_ net812 _01535_ net808 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08057__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09163_ _04212_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06375_ top.lcd.cnt_500hz\[8\] _01449_ _01495_ top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a311o_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08114_ _03230_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07804__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09094_ _04135_ _04138_ _04139_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ top.DUT.register\[13\]\[23\] net676 net651 top.DUT.register\[17\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a22o_1
XANTENNA__10781__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold920 top.DUT.register\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold931 top.DUT.register\[19\]\[8\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 top.DUT.register\[5\]\[28\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 top.DUT.register\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 top.DUT.register\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _01551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 top.DUT.register\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 top.DUT.register\[12\]\[10\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 top.DUT.register\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ net199 top.DUT.register\[2\]\[16\] net450 vssd1 vssd1 vccd1 vccd1 _00170_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07943__X _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net473 _04030_ _04034_ net394 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a22o_1
XANTENNA__06791__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ net271 _03811_ _03968_ net273 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o22a_1
XANTENNA__07335__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ top.DUT.register\[25\]\[28\] net637 net625 top.DUT.register\[16\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10021__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net2204 net174 net493 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07471__A_N _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ net188 net1741 net370 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10956__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08493__Y _03602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__A top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12510_ clknet_leaf_43_clk _00056_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13490_ clknet_leaf_107_clk _01036_ net952 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ clknet_leaf_53_clk top.ru.next_FetchedInstr\[4\] net1077 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08048__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09245__C1 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09796__B1 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ _06150_ net814 _06149_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__and3b_1
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11323_ net906 _05182_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10691__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ net909 _05012_ net403 net1237 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ net194 net2116 net439 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11185_ _04675_ net868 vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ net193 net2044 net442 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__mux2_1
XANTENNA_input39_X net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ net196 net2057 net447 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08397__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ clknet_leaf_59_clk _01351_ net1103 vssd1 vssd1 vccd1 vccd1 top.pad.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13757_ clknet_leaf_65_clk _01282_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10866__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ net2240 net190 net482 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12708_ clknet_leaf_30_clk _00254_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07964__A_N _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ clknet_leaf_79_clk _00010_ net1088 vssd1 vssd1 vccd1 vccd1 top.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ clknet_leaf_32_clk _00185_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 top.ramaddr\[9\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10454__X _04988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold216 top.DUT.register\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 top.DUT.register\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold238 top.DUT.register\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__S _04078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 top.DUT.register\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_4
X_09850_ _04843_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__nand2_1
XANTENNA__10106__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout718 _01559_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_4
Xfanout729 _01544_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07565__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ _03368_ _03882_ _03895_ net465 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o22ai_1
X_06993_ net324 _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and2_1
X_09781_ _01595_ _04198_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nor2_1
XANTENNA__06773__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ net398 _03154_ _03158_ net459 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07317__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _02522_ _03616_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nor2_1
XFILLER_0_205_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout173_A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__B top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07614_ top.DUT.register\[13\]\[11\] net676 net541 top.DUT.register\[5\]\[11\] _02730_
+ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a221o_1
X_08594_ _02666_ _03697_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_68_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ _02264_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10776__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout438_A _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07476_ top.DUT.register\[21\]\[7\] net571 net674 top.DUT.register\[19\]\[7\] _02592_
+ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06555__A top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _04260_ _04263_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11180__B net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06427_ net812 _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__nor2_2
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06274__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09778__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _04177_ _04198_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__or2_1
X_06358_ top.a1.instruction\[0\] top.a1.instruction\[1\] vssd1 vssd1 vccd1 vccd1 _01481_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ _03929_ _03946_ _03971_ _03991_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__or4_1
X_06289_ net1429 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[15\] sky130_fd_sc_hd__and2_1
XFILLER_0_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08028_ top.DUT.register\[6\]\[19\] net576 net544 top.DUT.register\[24\]\[19\] _03144_
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold750 top.DUT.register\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 top.DUT.register\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 top.DUT.register\[14\]\[13\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 top.DUT.register\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10016__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 top.DUT.register\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07556__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net615 _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__nand2_8
XFILLER_0_207_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12990_ clknet_leaf_37_clk _00536_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _05800_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__nand2_1
X_11872_ _05702_ net127 _05696_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ clknet_leaf_78_clk _01152_ net1085 vssd1 vssd1 vccd1 vccd1 top.ramload\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10823_ net1443 net249 net496 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
XANTENNA__10686__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06736__Y _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ clknet_leaf_47_clk _01088_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10754_ net258 net1904 net372 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XANTENNA__08009__X _03126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ clknet_leaf_41_clk _01019_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09218__C1 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ _04183_ net616 _04964_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09769__B1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ clknet_leaf_78_clk top.ru.next_FetchedData\[19\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ net1989 _06137_ net814 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07795__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ top.a1.row1\[2\] _05154_ _05161_ top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1
+ _05175_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12286_ net1190 _06096_ net1117 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ net871 _05109_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ net59 net884 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06755__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ net261 net2223 net445 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
X_11099_ net81 net878 net846 net1178 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22o_1
XANTENNA__11265__B top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07180__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ clknet_leaf_67_clk _01334_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10596__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _02440_ _02442_ _02444_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or4_4
XFILLER_0_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07261_ top.DUT.register\[22\]\[3\] net607 net729 top.DUT.register\[10\]\[3\] _02377_
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09000_ net1288 net890 _01797_ net622 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__a22o_1
X_06212_ net1361 _01428_ _01430_ _01385_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a22o_1
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_154_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07192_ top.DUT.register\[29\]\[10\] net784 net719 top.DUT.register\[26\]\[10\] _02308_
+ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08983__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_187_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _04891_ _04890_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 _04991_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_4
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_6
XANTENNA__07538__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout526 net528 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_8
X_09833_ net818 _04437_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__nor2_1
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_4
Xfanout559 _01677_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06746__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Right_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__B _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net820 _04299_ net817 top.pc\[8\] vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a2bb2o_1
X_06976_ top.DUT.register\[18\]\[20\] net779 net715 top.DUT.register\[9\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08715_ net306 _03423_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__nor2_1
X_09695_ top.a1.halfData\[1\] _01480_ _04710_ _04713_ net1102 vssd1 vssd1 vccd1 vccd1
+ _00117_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout555_A _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ _03743_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__or2_1
XANTENNA__07171__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ net302 _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__or2_1
XANTENNA__09448__C1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout722_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06556__Y _01673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07528_ top.DUT.register\[7\]\[13\] net572 net675 top.DUT.register\[13\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ _02569_ _02571_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__or3_1
XFILLER_0_146_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13834__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ net204 net1784 net507 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ net912 _01552_ _01597_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07777__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _05992_ _06000_ _05994_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_94_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13619__Q net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ _05876_ _05925_ _05929_ _05931_ _05927_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__o221ai_2
Xhold580 top.DUT.register\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 top.DUT.register\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ net864 _05035_ _05036_ net870 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1
+ _05037_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_125_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Left_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12973_ clknet_leaf_113_clk _00519_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11924_ _05777_ _05780_ _05781_ _05782_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__or4_4
XFILLER_0_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07162__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11855_ _05708_ _05713_ _05714_ _05707_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__and4b_1
X_10806_ net179 net1722 net411 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__mux2_1
XANTENNA__06195__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11786_ _05640_ _05645_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ clknet_leaf_98_clk _01071_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ net193 top.DUT.register\[24\]\[18\] net415 vssd1 vssd1 vccd1 vccd1 _00876_
+ sky130_fd_sc_hd__mux2_1
X_13456_ clknet_leaf_117_clk _01002_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10668_ net205 net1716 net420 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12407_ clknet_leaf_55_clk top.ru.next_FetchedData\[2\] net1097 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_max_cap353_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ clknet_leaf_5_clk _00933_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10599_ net218 net2267 net422 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07768__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08965__B2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12338_ top.pad.count\[0\] net920 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nand2_1
XANTENNA__06976__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ net1175 _06073_ _06087_ net1117 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08717__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__B2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06830_ top.DUT.register\[28\]\[27\] net739 net588 top.DUT.register\[20\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06761_ _01874_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nor2_2
X_08500_ _03377_ _03569_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a21o_1
X_09480_ _02089_ _04511_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__xnor2_1
X_06692_ _01808_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__inv_2
XFILLER_0_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07153__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06657__X _01774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ net303 _03541_ _03529_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06376__Y top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ _03402_ _03471_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07313_ top.DUT.register\[8\]\[7\] net595 net717 top.DUT.register\[9\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06536__C top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08293_ net285 _02428_ _03282_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_A _04208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ top.DUT.register\[28\]\[8\] net740 net762 top.DUT.register\[30\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ top.DUT.register\[27\]\[11\] net771 net759 top.DUT.register\[2\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout303_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__RESET_B net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout301 _01856_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_167_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout312 _01830_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
Xfanout323 net326 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
XANTENNA__08112__X _03229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__B _02028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 _01940_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
X_09816_ net203 net2218 net392 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
Xfanout378 net381 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
Xfanout389 _04969_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07931__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _03521_ net456 net535 _04755_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__o211a_4
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ top.DUT.register\[22\]\[21\] net605 net781 top.DUT.register\[1\]\[21\] _02075_
+ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout937_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11914__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ top.pad.keyCode\[5\] top.pad.keyCode\[4\] top.pad.keyCode\[7\] top.pad.keyCode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07144__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06567__X _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08629_ _02662_ _02821_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ _05466_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__xor2_2
XFILLER_0_166_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07447__A1 top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10964__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ _05414_ _05426_ _05431_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10817__X _04999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13310_ clknet_leaf_40_clk _00856_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07998__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ net262 net2249 net428 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13241_ clknet_leaf_58_clk _00787_ net1100 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ net2215 net140 net511 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__B2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ net1408 _04941_ net430 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__mux2_1
X_13172_ clknet_leaf_103_clk _00718_ net985 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06958__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _05969_ _05982_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _05886_ _05911_ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07574__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__X _04171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ top.a1.halfData\[2\] _05005_ _05023_ net864 vssd1 vssd1 vccd1 vccd1 _05024_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10204__S net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07383__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07922__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_4
XANTENNA__09014__A1_N _02714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12956_ clknet_leaf_16_clk _00502_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06477__X _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07135__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11907_ _05727_ _05762_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__xnor2_2
X_12887_ clknet_leaf_114_clk _00433_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _05697_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__or2_1
XANTENNA__09029__A1_N _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10874__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _05618_ _05620_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ clknet_leaf_29_clk _01054_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_151_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13439_ clknet_leaf_31_clk _00985_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08980_ net463 _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__nand2_1
X_07931_ top.DUT.register\[19\]\[25\] net674 net626 top.DUT.register\[16\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a22o_1
XANTENNA_wire359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _01981_ _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__or2_1
XANTENNA__07374__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _04608_ _04625_ _04626_ net823 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a31o_1
X_06813_ _01923_ _01925_ _01927_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07793_ top.DUT.register\[3\]\[29\] net691 net540 top.DUT.register\[5\]\[29\] _02909_
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09532_ _04560_ _04561_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06744_ top.DUT.register\[10\]\[28\] net728 net762 top.DUT.register\[30\]\[28\] _01860_
+ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a221o_1
XFILLER_0_195_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06675_ top.DUT.register\[5\]\[1\] net542 net630 top.DUT.register\[29\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a22o_1
X_09463_ _04475_ _04478_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_195_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ net291 _03384_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09394_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08345_ net284 _03375_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout420_A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout518_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ net284 _02070_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__nor2_1
XANTENNA__07659__A _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06652__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ top.DUT.register\[28\]\[9\] net740 net806 top.DUT.register\[15\]\[9\] _02343_
+ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a221o_1
XANTENNA__08929__A1 _03364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07158_ top.DUT.register\[19\]\[12\] net750 net748 top.DUT.register\[1\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07089_ top.DUT.register\[23\]\[15\] net732 net713 top.DUT.register\[25\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1111 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_2
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout131 net134 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
Xfanout142 _04957_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout153 _04932_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10024__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07365__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout175 _04878_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_1
XANTENNA__07904__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 _04858_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_137_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10959__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12810_ clknet_leaf_117_clk _00356_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13790_ clknet_leaf_70_clk _01315_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07117__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12741_ clknet_leaf_46_clk _00287_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12672_ clknet_leaf_15_clk _00218_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11623_ _05449_ _05450_ net207 vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__and3_1
XANTENNA__06891__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10694__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _05399_ _05380_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_146_Left_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10505_ net195 net2157 net379 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
XANTENNA__06643__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ _05342_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ clknet_leaf_26_clk _00770_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ net1311 net209 net509 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__mux2_1
XANTENNA__06760__X _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13552__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13155_ clknet_leaf_34_clk _00701_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10367_ net1540 net217 net430 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
X_12106_ _05897_ _05964_ _05957_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_209_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13086_ clknet_leaf_39_clk _00632_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10298_ net2191 net224 net521 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_89_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12037_ top.a1.dataIn\[4\] _05895_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_155_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07356__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10869__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07108__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ clknet_leaf_4_clk _00485_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06460_ top.DUT.register\[4\]\[0\] net581 net757 top.DUT.register\[3\]\[0\] _01576_
+ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08863__A _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06391_ top.pad.button_control.r_counter\[1\] top.pad.button_control.r_counter\[4\]
+ top.pad.button_control.r_counter\[3\] _01502_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__or4_1
XANTENNA__06882__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_164_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08130_ top.DUT.register\[6\]\[16\] net576 net675 top.DUT.register\[13\]\[16\] _03246_
+ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ net825 _03177_ _02617_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a21o_1
XANTENNA__10109__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07012_ _02122_ _02124_ _02126_ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07595__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net306 _03726_ _03886_ net269 _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_173_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07914_ _02023_ _03029_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__and2_1
X_08894_ _03941_ _03983_ net317 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07347__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ top.DUT.register\[23\]\[26\] net565 net557 top.DUT.register\[8\]\[26\] _02961_
+ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout370_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07776_ top.DUT.register\[18\]\[30\] net661 net646 top.DUT.register\[10\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ net133 _04534_ _04535_ _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o31a_1
X_06727_ top.DUT.register\[1\]\[3\] net706 net633 top.DUT.register\[27\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout635_A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09446_ net135 _04474_ _04480_ _04481_ net916 vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_182_Left_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06658_ net829 _01773_ _01754_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06873__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ top.pc\[15\] _04398_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06589_ top.DUT.register\[29\]\[0\] net628 net624 top.DUT.register\[16\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ _02845_ _03408_ _02555_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__o21a_1
XANTENNA__12693__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10019__S net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ net325 _01941_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11270_ net901 _05130_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_115_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10221_ net240 net1746 net383 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
XANTENNA__06740__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ net2272 net262 net527 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
XANTENNA__07050__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08013__A _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__A1 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ net614 _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__nand2_1
XANTENNA__07338__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 top.a1.dataInTemp\[7\] vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13481__RESET_B net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_42_clk _01365_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13773_ clknet_leaf_62_clk _01298_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_10985_ top.a1.halfData\[5\] _01433_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12724_ clknet_leaf_99_clk _00270_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ clknet_leaf_25_clk _00201_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11606_ _01396_ net207 _05437_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12586_ clknet_leaf_118_clk _00132_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _05334_ _05396_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold409 top.DUT.register\[18\]\[4\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06490__X _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06931__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _05323_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08369__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ clknet_leaf_111_clk _00753_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ net1587 net139 net515 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XANTENNA__07746__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _05252_ top.a1.dataIn\[29\] vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13138_ clknet_leaf_106_clk _00684_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07041__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13069_ clknet_leaf_114_clk _00615_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1109 top.DUT.register\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11125__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07762__A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ net400 _02589_ _02746_ _01615_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_179_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07561_ top.DUT.register\[2\]\[9\] net685 net677 top.DUT.register\[13\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09300_ net854 _01635_ net619 vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__o21a_1
X_06512_ _01598_ _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__nand2_1
X_07492_ _02602_ _02604_ _02606_ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12472__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _04277_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__or2_1
XANTENNA__06855__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06443_ top.a1.instruction\[15\] top.a1.instruction\[16\] net810 _01542_ vssd1 vssd1
+ vccd1 vccd1 _01560_ sky130_fd_sc_hd__and4_4
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06374_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__or4_1
X_09162_ _04213_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08113_ _02068_ _03228_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_211_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09093_ _03813_ _03828_ _04140_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__or4b_1
XFILLER_0_43_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ top.DUT.register\[22\]\[23\] net552 net639 top.DUT.register\[9\]\[23\] _03160_
+ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07937__A _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07280__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold910 top.DUT.register\[17\]\[7\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 top.DUT.register\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold932 top.DUT.register\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 top.DUT.register\[6\]\[30\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 top.DUT.register\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold965 top.DUT.register\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 top.DUT.register\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09106__D_N _03229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold987 top.DUT.register\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold998 top.DUT.register\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net205 net1661 net452 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout585_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net306 _03707_ _03571_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _03885_ _03967_ net291 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10302__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ top.DUT.register\[3\]\[28\] net692 net562 top.DUT.register\[20\]\[28\] _02944_
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_86_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06288__A top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_190_Left_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _02869_ _02871_ _02873_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07099__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ net192 net2259 net370 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
XANTENNA__06575__X _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09429_ net135 _04458_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06846__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ clknet_leaf_54_clk top.ru.next_FetchedInstr\[3\] net1076 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09886__X _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12371_ top.pad.button_control.r_counter\[10\] top.pad.button_control.r_counter\[9\]
+ _06146_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__and3_1
XANTENNA__10972__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09796__B2 top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _05183_ _05188_ _05189_ _05187_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__or4b_1
XANTENNA__07271__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11253_ _05126_ net1246 net402 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07559__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net198 net1545 net438 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
XANTENNA__07023__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _01441_ _01444_ _05092_ top.busy_o vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__o22a_1
XFILLER_0_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10135_ net196 net2086 net443 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__B _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ net199 top.DUT.register\[4\]\[16\] net446 vssd1 vssd1 vccd1 vccd1 _00234_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10212__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13825_ clknet_leaf_71_clk _01350_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13756_ clknet_leaf_65_clk _01281_ net1099 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10968_ net1474 net193 net481 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XANTENNA__09484__B1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12707_ clknet_leaf_34_clk _00253_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12544__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09302__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06837__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13687_ clknet_leaf_74_clk _01227_ net1089 vssd1 vssd1 vccd1 vccd1 top.busy_o sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ net2231 net203 net407 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
X_12638_ clknet_leaf_37_clk _00184_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10882__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ clknet_leaf_62_clk _00115_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07262__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 top.DUT.register\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold217 top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 top.DUT.register\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06470__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 top.DUT.register\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout708 net710 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_8
Xfanout719 _01548_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
XANTENNA__13332__RESET_B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08800_ _03232_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07763__Y _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ top.pc\[12\] _04198_ _04359_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ _02099_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__nor2_2
XANTENNA__07970__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ net475 _03153_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09172__C1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ net398 _03254_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nor2_1
XANTENNA__10122__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06525__A1 top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07613_ top.DUT.register\[1\]\[11\] net704 net557 top.DUT.register\[8\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ _03671_ _02823_ _02820_ _02284_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a2bb2o_1
X_07544_ net829 net333 net468 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09212__A _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06828__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ top.DUT.register\[14\]\[7\] net665 net658 top.DUT.register\[28\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1075_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__B top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _04260_ _04263_ net822 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__a21oi_1
X_06426_ _01527_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__A1 _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _02519_ _04197_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__nand2_2
X_06357_ _01480_ vssd1 vssd1 vccd1 vccd1 top.edg2.button_i sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10792__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09076_ net296 net279 _03460_ _04051_ _02517_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__a311o_1
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06288_ top.ramload\[14\] net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08158__C_N _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08027_ top.DUT.register\[31\]\[19\] net667 net639 top.DUT.register\[9\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold740 top.DUT.register\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06290__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold751 top.DUT.register\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold762 top.DUT.register\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 top.DUT.register\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 top.DUT.register\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 top.a1.row2\[41\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _04729_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__nor2_2
X_08929_ _03364_ _04013_ _04014_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11940_ _05787_ _05797_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__nand2_1
XANTENNA__10032__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11871_ _05696_ _05702_ net127 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__and3_1
XANTENNA__10967__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ clknet_leaf_74_clk _01151_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramload\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ net1993 net253 net495 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13541_ clknet_leaf_47_clk _01087_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ net261 net2102 net373 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06819__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13472_ clknet_leaf_12_clk _01018_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10684_ net141 net1728 net421 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09769__A1 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ clknet_leaf_74_clk top.ru.next_FetchedData\[18\] net1086 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12354_ top.pad.button_control.r_counter\[4\] top.pad.button_control.r_counter\[3\]
+ _06135_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__and3_1
XANTENNA__07244__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06481__A top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11305_ top.a1.row1\[18\] _05155_ _05160_ top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1
+ _05174_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12285_ _06096_ _06097_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10207__S net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11328__B2 top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _05118_ net1323 net402 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06536__A_N top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08907__A_N _03995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ net924 net1268 net876 _05083_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a31o_1
XANTENNA__07952__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ net243 net1656 net443 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__mux2_1
X_11098_ net80 net879 net847 net1171 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11265__C top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10049_ net614 _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12725__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10877__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13808_ clknet_leaf_68_clk _01333_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ clknet_leaf_68_clk _00004_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07260_ top.DUT.register\[23\]\[3\] net732 _01546_ top.DUT.register\[16\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08680__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06211_ _01425_ _00017_ _01420_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__and3b_1
XFILLER_0_170_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07191_ top.DUT.register\[13\]\[10\] net788 net715 top.DUT.register\[9\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_154_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08432__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08983__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06994__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ top.pc\[24\] _04557_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09906__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _04988_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_8
Xfanout516 _04985_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_6
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_6
XANTENNA__07493__Y _02610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _04824_ _04827_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout549 _01687_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_206_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_206_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _02519_ _04197_ _04767_ net457 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a31o_2
X_06975_ top.DUT.register\[21\]\[20\] net608 net734 top.DUT.register\[12\]\[20\] _02091_
+ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout283_A _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ net270 _03635_ _03811_ net277 _03812_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a221oi_2
X_09694_ _04700_ _04704_ _04711_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__or4_1
XFILLER_0_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08645_ _03361_ _03459_ net307 vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout450_A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10787__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08576_ _03594_ _03680_ net289 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07527_ top.DUT.register\[2\]\[13\] net683 net540 top.DUT.register\[5\]\[13\] _02643_
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout715_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ top.DUT.register\[4\]\[6\] net551 _02572_ _02574_ vssd1 vssd1 vccd1 vccd1
+ _02575_ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06409_ net809 _01525_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__nor2_1
XANTENNA__06572__Y _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07389_ top.DUT.register\[10\]\[4\] net728 net772 top.DUT.register\[27\]\[4\] _02505_
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09128_ top.a1.instruction\[9\] top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ _04181_ sky130_fd_sc_hd__and2_1
XANTENNA__08423__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07226__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10027__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ _04015_ _04037_ _04058_ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09816__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ _05898_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and2_1
Xhold570 top.DUT.register\[30\]\[1\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 top.DUT.register\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 top.DUT.register\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ top.a1.data\[2\] net796 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__or2_1
XANTENNA__09923__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ clknet_leaf_115_clk _00518_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _05780_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nor2_1
XANTENNA__10697__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11854_ _05713_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10805_ net186 net1870 net410 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ _05643_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13659__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13524_ clknet_leaf_97_clk _01070_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10736_ net198 net1713 net415 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07465__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13455_ clknet_leaf_20_clk _01001_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ net209 net1621 net418 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06482__Y _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ clknet_leaf_54_clk top.ru.next_FetchedData\[1\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07217__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_118_clk _00932_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10598_ net222 net2265 net423 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__mux2_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__clkbuf_4
X_12337_ top.lcd.cnt_500hz\[14\] _06127_ _06128_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12268_ _06074_ _06079_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nand2_1
XANTENNA__08717__A2 _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ net1269 net405 net369 _05110_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a22o_1
X_12199_ _06051_ _06056_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__xor2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07925__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire349_A _02283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06760_ _01863_ _01864_ _01865_ _01876_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__or4_4
X_06691_ top.a1.instruction\[25\] net857 _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_201_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ net281 _03532_ _03531_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_65_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10400__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ net308 _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08102__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07312_ net297 _02428_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07456__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06664__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07243_ top.DUT.register\[3\]\[8\] net783 net724 top.DUT.register\[16\]\[8\] _02359_
+ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06325__S _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ top.DUT.register\[11\]\[11\] net767 net589 top.DUT.register\[20\]\[11\] _02290_
+ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a221o_1
XANTENNA__08405__B2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1038_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 _01856_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout498_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_7__f_clk_X clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07664__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_2
XANTENNA__07916__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09815_ _03758_ net455 net534 _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__o211a_4
XFILLER_0_185_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout379 net381 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_4
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout665_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ top.pc\[5\] net817 net457 _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a211o_1
X_06958_ top.DUT.register\[4\]\[21\] net582 net708 top.DUT.register\[7\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07680__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _04694_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ top.DUT.register\[21\]\[24\] net610 net587 top.DUT.register\[24\]\[24\] _02005_
+ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout832_A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ net394 _03721_ _03727_ net474 _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__a221o_1
XANTENNA__10310__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07695__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ net281 _03439_ _03572_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_59_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08644__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__nand2_1
XANTENNA__08644__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13435__RESET_B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ net242 net1640 net427 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ clknet_leaf_37_clk _00786_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10452_ net1415 net143 net511 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__mux2_1
XANTENNA__13857__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ clknet_leaf_107_clk _00717_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ net1609 net150 net431 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ _05977_ _05980_ _05970_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12053_ _05894_ _05913_ _05884_ _05886_ _05890_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07907__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ top.a1.dataInTemp\[2\] net798 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__or2_1
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout891 _01438_ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_12955_ clknet_leaf_0_clk _00501_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ _05763_ _05766_ _05764_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07686__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ clknet_leaf_14_clk _00432_ net986 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ top.a1.dataIn\[7\] _05682_ _05686_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__and3_1
XANTENNA__06894__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08635__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11768_ _05626_ _05627_ _05622_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ clknet_leaf_34_clk _01053_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10719_ net243 net1644 net415 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
X_11699_ _05559_ _05523_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_151_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13438_ clknet_leaf_38_clk _00984_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10890__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ clknet_leaf_57_clk _00915_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_184_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07071__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11287__A top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ top.DUT.register\[13\]\[25\] net678 net665 top.DUT.register\[14\]\[25\] _03046_
+ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07861_ net828 _02977_ _02618_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__o21a_1
XANTENNA__12740__RESET_B net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ _04608_ _04626_ _04625_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a21oi_1
X_06812_ top.DUT.register\[6\]\[31\] net599 net764 top.DUT.register\[19\]\[31\] _01928_
+ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a221o_1
X_07792_ top.DUT.register\[1\]\[29\] net703 net683 top.DUT.register\[2\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _04561_ _04560_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and2b_1
X_06743_ top.DUT.register\[23\]\[28\] net731 net724 top.DUT.register\[16\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10130__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _04495_ _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nand2_1
X_06674_ top.DUT.register\[6\]\[1\] net578 net567 top.DUT.register\[23\]\[1\] _01790_
+ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a221o_1
X_08413_ _02837_ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_195_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09393_ top.pc\[15\] _04398_ top.pc\[16\] vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ net463 _03443_ _03452_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__a211o_1
XANTENNA__07429__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ net270 _03386_ _03389_ net277 vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout413_A _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07226_ top.DUT.register\[29\]\[9\] net786 net751 top.DUT.register\[19\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07157_ top.DUT.register\[6\]\[12\] net596 net804 top.DUT.register\[15\]\[12\] _02269_
+ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07062__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07088_ top.DUT.register\[14\]\[15\] net794 net582 top.DUT.register\[4\]\[15\] _02204_
+ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout782_A _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1110 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10305__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_4_1__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout132 net134 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09890__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 net146 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
Xfanout154 _04923_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _04905_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_199_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout176 _04878_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 net190 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _04833_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_202_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09729_ net242 net2216 net391 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ clknet_leaf_31_clk _00286_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11363__C top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08793__X _03888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13616__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12671_ clknet_leaf_23_clk _00217_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08953__B _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ _05446_ _05475_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _05404_ _05407_ _05409_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08093__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ net200 net1740 net378 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__mux2_1
X_11484_ _05269_ _05306_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ clknet_leaf_56_clk _00769_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10435_ net1430 net214 net510 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ clknet_leaf_11_clk _00700_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ net1310 net219 net431 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12105_ top.a1.dataIn\[3\] _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__nor2_1
XANTENNA__06800__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ clknet_leaf_120_clk _00631_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10215__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10297_ net1915 net230 net523 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
X_12036_ top.a1.dataIn\[4\] _05895_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11273__C top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ clknet_leaf_116_clk _00484_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12439__Q top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10885__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ clknet_leaf_40_clk _00415_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08863__B _03954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06390_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[8\]
+ top.pad.button_control.r_counter\[6\] top.pad.button_control.r_counter\[2\] vssd1
+ vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__or4_1
XFILLER_0_173_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09805__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ _03161_ _03163_ _03167_ _03176_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__or4_2
XANTENNA__07831__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ top.DUT.register\[5\]\[19\] net601 net588 top.DUT.register\[20\]\[19\] _02127_
+ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07044__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__A _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10125__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ net293 _03967_ _04048_ net279 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_164_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07913_ _02023_ _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nor2_1
X_08893_ net325 _01981_ _03344_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ top.DUT.register\[3\]\[26\] net692 net669 top.DUT.register\[31\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a22o_1
XANTENNA__07898__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07775_ top.DUT.register\[8\]\[30\] net559 net634 top.DUT.register\[27\]\[30\] _02891_
+ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ net136 _04540_ _04545_ net822 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__o22a_1
X_06726_ _01836_ _01838_ _01840_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__or4_1
XFILLER_0_189_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08847__B2 _02024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13098__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09445_ _04475_ _04478_ _04479_ net821 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10795__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06657_ net828 _01773_ _01754_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout530_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _04414_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06588_ _01672_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08327_ net309 _03440_ _03433_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09272__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07283__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _03282_ _03366_ net463 _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__a31o_1
XANTENNA__07822__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09100__D _03054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07209_ _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__inv_2
XANTENNA__09024__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ _03303_ _03304_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10220_ net614 _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ net1526 net243 net526 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XANTENNA__10035__S net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09028__A1_N _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10082_ _04732_ _04965_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nor2_1
X_13841_ clknet_leaf_42_clk _01364_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06561__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13772_ clknet_leaf_73_clk _01297_ net1120 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net869 net864 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06849__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ clknet_leaf_108_clk _00269_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ clknet_leaf_96_clk _00200_ net1000 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11605_ _01396_ net207 vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12585_ clknet_leaf_8_clk _00131_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07274__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ _05337_ _05366_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__xnor2_1
Xwire341 _02407_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_2
Xwire352 _02194_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11467_ _05281_ _05283_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07026__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ clknet_leaf_104_clk _00752_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ net1506 net143 net516 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11398_ _05246_ _05247_ _05252_ _05253_ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ clknet_leaf_7_clk _00683_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10349_ net2022 net156 net517 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ clknet_leaf_2_clk _00614_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05876_ _05878_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nand2_1
XANTENNA_wire331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ top.DUT.register\[17\]\[9\] net653 _02674_ _02676_ vssd1 vssd1 vccd1 vccd1
+ _02677_ sky130_fd_sc_hd__a211o_1
X_06511_ _01620_ _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__or2_1
X_07491_ top.DUT.register\[20\]\[7\] net562 net633 top.DUT.register\[27\]\[7\] _02607_
+ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09230_ top.pc\[6\] _04254_ top.pc\[7\] vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06442_ net811 _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__nor2_4
XFILLER_0_29_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09161_ _01753_ net341 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__and2_1
XANTENNA__08057__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06373_ net34 top.ru.state\[0\] _01492_ vssd1 vssd1 vccd1 vccd1 top.ru.next_read_i
+ sky130_fd_sc_hd__and3_1
X_08112_ _02068_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__or2_2
XANTENNA__07265__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__B2 top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09092_ _03597_ _03614_ _04141_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_211_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07804__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08043_ top.DUT.register\[21\]\[23\] net569 net560 top.DUT.register\[20\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a22o_1
Xhold900 top.DUT.register\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09006__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold911 top.DUT.register\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 top.DUT.register\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold933 top.DUT.register\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold944 top.DUT.register\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08114__A _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold955 top.DUT.register\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 top.DUT.register\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 top.DUT.register\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net208 net1764 net450 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
Xhold988 top.DUT.register\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold999 top.DUT.register\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06240__B2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ net279 net470 _03503_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_110_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06791__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout578_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _03923_ _03966_ net318 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07827_ top.DUT.register\[24\]\[28\] net546 net661 top.DUT.register\[18\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a22o_1
XANTENNA__06288__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07758_ top.DUT.register\[6\]\[31\] net579 net574 top.DUT.register\[7\]\[31\] _02874_
+ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06709_ top.DUT.register\[30\]\[4\] net697 net562 top.DUT.register\[20\]\[4\] _01825_
+ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a221o_1
X_07689_ top.DUT.register\[24\]\[12\] net544 _02805_ vssd1 vssd1 vccd1 vccd1 _02806_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ net131 _04453_ _04463_ _04464_ net916 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o221a_1
XFILLER_0_192_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ _04398_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08048__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09245__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11052__A1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12370_ top.pad.button_control.r_counter\[9\] _06146_ top.pad.button_control.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ net900 _05184_ _05165_ _05151_ _05140_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07008__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net871 _05113_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__and2_1
XANTENNA__13638__Q net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ net199 top.DUT.register\[8\]\[16\] net438 vssd1 vssd1 vccd1 vccd1 _00362_
+ sky130_fd_sc_hd__mux2_1
X_11183_ wb.curr_state\[0\] net877 _01443_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ net202 net2018 net442 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__mux2_1
XANTENNA__11107__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10065_ net203 net2297 net448 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XANTENNA__06479__A top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13824_ clknet_leaf_70_clk _01349_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ clknet_leaf_65_clk _01280_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10967_ net1496 net195 net481 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09302__B _04345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ clknet_leaf_11_clk _00252_ net974 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10898_ net1670 net210 net406 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
X_13686_ clknet_leaf_77_clk _01226_ net1081 vssd1 vssd1 vccd1 vccd1 top.pc\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ clknet_leaf_120_clk _00183_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09729__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ clknet_leaf_62_clk _00114_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08995__B1 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ _05372_ _05375_ _05379_ _05377_ _05363_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__a32o_1
X_12499_ clknet_leaf_87_clk _00046_ net1018 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold207 top.ramaddr\[23\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 top.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 top.DUT.register\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12452__Q top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_6
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06991_ _02101_ _02103_ _02105_ _02107_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__or4_2
XANTENNA__06773__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net271 _03661_ _03826_ net274 _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o221a_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10403__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ net312 _02201_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07612_ _02722_ _02724_ _02726_ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__or4_1
X_08592_ net1536 net858 net836 _03696_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
X_07543_ _02644_ _02646_ _02650_ _02659_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__nor4_1
XFILLER_0_88_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout159_A _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07474_ top.a1.instruction\[28\] net857 _01615_ _02590_ vssd1 vssd1 vccd1 vccd1 _02591_
+ sky130_fd_sc_hd__a22oi_4
X_09213_ _04261_ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nand2_1
X_06425_ top.a1.instruction\[17\] top.a1.instruction\[18\] net830 vssd1 vssd1 vccd1
+ vccd1 _01542_ sky130_fd_sc_hd__and3b_1
XANTENNA__09227__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09227__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1068_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07238__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _04179_ _04180_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__o21ba_1
X_06356_ top.pad.button_control.debounce_dly top.pad.button_control.debounce vssd1
+ vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__and2b_2
XANTENNA__12231__B1 _05094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09075_ _04124_ _04125_ _04126_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__or4_1
X_06287_ net1180 net897 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ top.DUT.register\[11\]\[19\] net699 net696 top.DUT.register\[30\]\[19\] _03142_
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold730 top.DUT.register\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 top.DUT.register\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold752 top.a1.row2\[16\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 top.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold774 top.DUT.register\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 top.DUT.register\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 top.DUT.register\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout862_A _05053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ top.a1.instruction\[7\] top.a1.instruction\[8\] net744 vssd1 vssd1 vccd1
+ vccd1 _04959_ sky130_fd_sc_hd__nand3b_2
XANTENNA__06764__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net473 _04007_ _04010_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09106__C _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ net473 _03945_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__nand2_1
XANTENNA__06586__X _01703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ net1369 net265 net496 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09466__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13540_ clknet_leaf_31_clk _01086_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10752_ net240 net1798 net371 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XANTENNA__07477__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ clknet_leaf_23_clk _01017_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ net145 net2007 net421 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09218__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ clknet_leaf_79_clk top.ru.next_FetchedData\[17\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_164_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__A2 _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08977__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12353_ _06137_ _06138_ net814 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11304_ net1207 net843 _05173_ net1115 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12284_ net1965 _06095_ net1117 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11235_ net871 _05026_ _05038_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09137__X _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ net58 net884 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net614 _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nand2_1
XANTENNA__10223__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ net79 net884 net849 net1155 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a22o_1
X_10048_ _04738_ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__nor2_1
Xhold90 top.ramstore\[27\] vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07180__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ clknet_leaf_69_clk _01332_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11999_ _05823_ _05827_ _05859_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09032__B _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13738_ clknet_leaf_67_clk _00003_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10893__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ clknet_leaf_90_clk _01210_ net1010 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06210_ net2065 _01428_ _01429_ net907 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ top.DUT.register\[15\]\[10\] net804 net800 top.DUT.register\[31\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09090__C1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08983__A3 _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06994__A2 _02089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09900_ top.pc\[23\] _02615_ _04882_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a21o_1
XANTENNA__10527__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout506 _04988_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_4
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout517 _04983_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_6
X_09831_ _04824_ _04827_ _04192_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_169_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout528 _04972_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_4
Xfanout539 _03291_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_4
XANTENNA__06746__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10133__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ top.DUT.register\[13\]\[20\] net788 net760 top.DUT.register\[30\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22o_1
XANTENNA__09207__B _01808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ net457 _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_206_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ net302 _03414_ net305 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o21a_1
X_09693_ _04692_ _04696_ _04703_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout276_A _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net476 _02717_ _02720_ net458 _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a221o_1
XANTENNA__07171__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ _03633_ _03679_ net314 vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07526_ top.DUT.register\[30\]\[13\] net695 net631 top.DUT.register\[27\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ top.DUT.register\[14\]\[6\] net665 net645 top.DUT.register\[10\]\[6\] _02573_
+ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09877__B _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06408_ _01389_ _01519_ _01523_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__or3_1
XFILLER_0_162_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08273__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07388_ top.DUT.register\[29\]\[4\] net786 net757 top.DUT.register\[3\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09127_ _01387_ _01490_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nor2_1
X_06339_ _01334_ _01330_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__and2b_1
XANTENNA__10308__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ _03953_ _03965_ _03994_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__and4_1
XFILLER_0_102_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _03116_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__or2_2
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold560 top.DUT.register\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold571 top.DUT.register\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ top.a1.dataInTemp\[6\] _05009_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__or2_1
Xhold582 top.DUT.register\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 top.DUT.register\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10043__S net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__B _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ clknet_leaf_6_clk _00517_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10978__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _05781_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__or2_1
XANTENNA__07698__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11853_ _05671_ _05689_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09439__A1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ net187 net2014 net410 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__mux2_1
X_11784_ _05607_ _05632_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08111__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ clknet_leaf_109_clk _01069_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ net200 net2190 net414 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XANTENNA__13260__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13454_ clknet_leaf_94_clk _01000_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10666_ net212 net2325 net418 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__mux2_1
XANTENNA__07870__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06492__A _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12405_ clknet_leaf_54_clk top.ru.next_FetchedData\[0\] net1096 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10218__S net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13385_ clknet_leaf_26_clk _00931_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10597_ net223 net2285 net422 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
X_12336_ top.lcd.cnt_500hz\[14\] _06127_ net743 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a21boi_1
XANTENNA__06976__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12267_ _06080_ _06086_ net1117 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__o21a_1
XANTENNA__08178__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output72_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ top.a1.dataInTemp\[8\] top.a1.data\[8\] net798 vssd1 vssd1 vccd1 vccd1 _05110_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09375__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12198_ top.a1.dataIn\[1\] _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or3_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__06728__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ net922 net1316 net874 _05074_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_182_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10888__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06690_ _01804_ _01803_ net401 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XANTENNA__07153__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06900__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ net301 _03472_ _03471_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07311_ _02418_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nor2_8
XFILLER_0_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ net308 _03405_ _03390_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_190_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07242_ top.DUT.register\[29\]\[8\] net786 net713 top.DUT.register\[25\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07173_ top.DUT.register\[12\]\[11\] net735 net750 top.DUT.register\[19\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a22o_1
XANTENNA__10128__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09917__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06967__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout303 net305 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
Xfanout314 net316 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13736__Q top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
XANTENNA_fanout393_A _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09814_ net816 _04811_ _04812_ _04807_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a31o_1
Xfanout369 _05108_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_2
XFILLER_0_185_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07392__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ net820 _04256_ top.a1.dataIn\[5\] net813 vssd1 vssd1 vccd1 vccd1 _04754_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout560_A _01673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ top.DUT.register\[27\]\[21\] net771 net585 top.DUT.register\[24\]\[21\] _02073_
+ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout658_A _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ top.pad.keyCode\[0\] top.pad.keyCode\[2\] top.pad.keyCode\[3\] top.pad.keyCode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or4b_1
XFILLER_0_179_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06888_ top.DUT.register\[26\]\[24\] net722 net595 top.DUT.register\[8\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
XANTENNA__07144__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ _02641_ net458 _03722_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08558_ net304 _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ top.DUT.register\[11\]\[14\] net699 net659 top.DUT.register\[18\]\[14\] _02625_
+ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ _03572_ _03588_ _03587_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ net616 _04960_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__nand2_1
XANTENNA__09400__B _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07852__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ net1360 net148 net509 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__mux2_1
XANTENNA__10038__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13475__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13170_ clknet_leaf_106_clk _00716_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07604__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ net1979 net156 net430 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ _05978_ _05980_ _05966_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06958__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ _05867_ _05872_ _05880_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__or4_1
Xhold390 top.DUT.register\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ top.a1.halfData\[2\] net796 vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__or2_1
Xfanout870 _04680_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_2
XANTENNA__07383__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout881 net883 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_1
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12500__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_19_clk _00500_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07135__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 top.DUT.register\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ _05752_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12885_ clknet_leaf_101_clk _00431_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08883__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__Y _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11836_ _05682_ _05686_ top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12650__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08096__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ _05626_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ clknet_leaf_11_clk _01052_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07843__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ net616 _04975_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2_1
X_11698_ _05517_ _05537_ _05538_ _05534_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_151_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13437_ clknet_leaf_119_clk _00983_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10649_ net149 net1717 net374 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08399__B2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__B1 _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13368_ clknet_leaf_33_clk _00914_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12319_ top.lcd.cnt_500hz\[7\] _06115_ top.lcd.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1
+ _06117_ sky130_fd_sc_hd__a21o_1
X_13299_ clknet_leaf_108_clk _00845_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11287__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _02967_ _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nor2_2
XANTENNA__07374__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ top.DUT.register\[23\]\[31\] net732 net774 top.DUT.register\[2\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a22o_1
X_07791_ top.DUT.register\[8\]\[29\] net556 net643 top.DUT.register\[10\]\[29\] _02907_
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a221o_1
X_06742_ net472 _01802_ net272 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or3_1
X_09530_ _04541_ _04542_ _04543_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10411__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09461_ _02099_ _02108_ _04494_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__or3_1
X_06673_ top.DUT.register\[24\]\[1\] net546 net649 top.DUT.register\[12\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a22o_1
XANTENNA__09979__Y _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _02550_ _03496_ _02588_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09392_ top.pc\[15\] top.pc\[16\] _04398_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_195_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08343_ net464 _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09823__A1 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout239_A _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__B2 top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _03387_ _03388_ net291 vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ top.DUT.register\[17\]\[9\] net753 _02330_ _02341_ vssd1 vssd1 vccd1 vccd1
+ _02342_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ top.DUT.register\[5\]\[12\] net600 net588 top.DUT.register\[20\]\[12\] _02272_
+ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07087_ top.DUT.register\[21\]\[15\] net610 net709 top.DUT.register\[7\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09890__B _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout155 _04923_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_1
XANTENNA__07365__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout166 net169 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08562__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__B2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _04878_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_199_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout188 net190 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout942_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ _03104_ _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__and2b_2
X_09728_ _03290_ net455 net534 _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o211a_2
XFILLER_0_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07117__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _04676_ net868 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11363__D top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12670_ clknet_leaf_40_clk _00216_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08078__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ _05443_ _05448_ net207 vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09814__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07825__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _05393_ _05411_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10503_ net206 net2315 net380 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
X_11483_ _05307_ _05308_ _05330_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ net1578 net216 net509 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
X_13222_ clknet_leaf_50_clk _00768_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ clknet_leaf_41_clk _00699_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10365_ net1497 net225 net430 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12104_ _05898_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__xnor2_4
X_13084_ clknet_leaf_81_clk _00630_ net1079 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10296_ net1406 net232 net523 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__mux2_1
X_12035_ _05892_ _05894_ top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08002__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12538__RESET_B net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06564__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10231__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__A1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07106__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12937_ clknet_leaf_8_clk _00483_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12868_ clknet_leaf_28_clk _00414_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_199_Right_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08069__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_177_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _05645_ _05678_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_32_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09805__A1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ clknet_leaf_32_clk _00345_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07816__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07292__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06951__Y _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07010_ top.DUT.register\[3\]\[19\] net756 net750 top.DUT.register\[19\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a22o_1
XANTENNA__07495__B _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10406__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07595__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ net294 _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ net828 _03028_ _02618_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__o21a_1
X_08892_ _03009_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__xor2_2
XANTENNA__07347__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__B1 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ top.DUT.register\[13\]\[26\] net676 net636 top.DUT.register\[25\]\[26\] _02959_
+ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_87_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout189_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ top.DUT.register\[2\]\[30\] net686 net642 top.DUT.register\[9\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07016__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09513_ _04541_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__xor2_1
X_06725_ top.DUT.register\[26\]\[3\] net682 net559 top.DUT.register\[8\]\[3\] _01841_
+ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout356_A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _04478_ _04479_ _04475_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a21oi_1
X_06656_ _01763_ _01772_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nor2_4
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _04408_ _04412_ _04413_ net821 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__a31o_1
X_06587_ top.a1.instruction\[22\] top.a1.instruction\[23\] net799 vssd1 vssd1 vccd1
+ vccd1 _01704_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout523_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08326_ net283 _03439_ _03437_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08257_ net472 net272 _03360_ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_201_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07208_ _02320_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__nor2_4
XFILLER_0_6_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08188_ net322 _02284_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07139_ top.DUT.register\[2\]\[13\] net758 net754 top.DUT.register\[18\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10316__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07586__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _04183_ net615 _04964_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ net139 net1674 net449 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
XANTENNA__09732__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_42_clk _01363_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10051__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13771_ clknet_leaf_73_clk _01296_ net1120 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_10983_ net908 top.a1.state\[0\] vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ clknet_leaf_106_clk _00268_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12653_ clknet_leaf_115_clk _00199_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11604_ _05456_ _05463_ _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08980__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12584_ clknet_leaf_25_clk _00130_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11535_ _05347_ _05350_ _05365_ _05391_ _05348_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a32o_2
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ _05325_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13205_ clknet_leaf_101_clk _00751_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ net1470 net147 net513 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
XANTENNA__10226__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11397_ top.a1.dataIn\[27\] _05255_ _05256_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_104_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13136_ clknet_leaf_117_clk _00682_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10348_ net1482 net161 net519 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XANTENNA__06785__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10279_ net168 net1559 net437 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__mux2_1
X_13067_ clknet_leaf_6_clk _00613_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07329__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11125__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _05868_ _05875_ _05877_ _05873_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_136_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10896__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06510_ _01497_ _01621_ _01622_ _01624_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__or4b_1
X_07490_ top.DUT.register\[1\]\[7\] net705 net550 top.DUT.register\[4\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06441_ _01518_ _01542_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _01753_ net341 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__nor2_1
X_06372_ _01494_ vssd1 vssd1 vccd1 vccd1 top.ru.next_write_i sky130_fd_sc_hd__inv_2
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08111_ net828 _03227_ net468 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09091_ _03510_ _04142_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08042_ _03082_ _03106_ _03132_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or4_1
Xhold901 top.DUT.register\[17\]\[28\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 top.DUT.register\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold923 top.DUT.register\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10136__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold934 top.DUT.register\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 top.DUT.register\[8\]\[27\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold956 top.DUT.register\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 top.DUT.register\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold978 top.DUT.register\[20\]\[2\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net212 net2320 net450 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__mux2_1
Xhold989 top.DUT.register\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06776__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ net477 _02927_ _02932_ net459 _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_95_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08517__B2 _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _01983_ _02004_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout473_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ top.DUT.register\[9\]\[28\] net640 net628 top.DUT.register\[29\]\[28\] _02942_
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07757_ top.DUT.register\[8\]\[31\] net558 net637 top.DUT.register\[25\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout640_A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06708_ top.DUT.register\[26\]\[4\] net682 net625 top.DUT.register\[16\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a22o_1
X_07688_ top.DUT.register\[18\]\[12\] net659 net631 top.DUT.register\[27\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a22o_1
X_09427_ _04461_ _04462_ net821 vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a21o_1
X_06639_ top.DUT.register\[7\]\[2\] net573 net652 top.DUT.register\[17\]\[2\] _01755_
+ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_A top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13837__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09358_ top.pc\[14\] _04368_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ net309 _03423_ _03390_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_23_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09289_ net915 top.pc\[10\] _04333_ net910 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__o211a_1
X_11320_ net900 _05127_ _05130_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11251_ _05125_ net1354 net402 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12883__RESET_B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net205 net1872 net440 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
X_11182_ net911 top.pc\[0\] _05089_ _05091_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a31o_1
XANTENNA__06767__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11666__A top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ net203 net1944 net444 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__mux2_1
XANTENNA__09407__Y _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ net208 net2344 net446 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_202_Right_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07192__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09423__X _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_70_clk _01348_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13754_ clknet_leaf_65_clk _01279_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08186__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ net1532 net201 net481 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12705_ clknet_leaf_41_clk _00251_ net1070 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13685_ clknet_leaf_67_clk _01225_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10897_ net1546 net214 net406 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ clknet_leaf_18_clk _00182_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07597__Y _02714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ clknet_leaf_62_clk _00113_ net1110 vssd1 vssd1 vccd1 vccd1 top.a1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_156_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08995__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11518_ _05361_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nor2_1
X_12498_ clknet_leaf_87_clk _00045_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold208 top.DUT.register\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold219 top.DUT.register\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06470__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11449_ top.a1.dataIn\[18\] _05243_ _05269_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06758__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10751__Y _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13119_ clknet_leaf_31_clk _00665_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ top.DUT.register\[16\]\[20\] net725 net589 top.DUT.register\[20\]\[20\] _02106_
+ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a221o_1
XANTENNA__07970__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ _03257_ _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07183__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ top.DUT.register\[21\]\[11\] net569 net684 top.DUT.register\[2\]\[11\] _02727_
+ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09012__A1_N _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08591_ net902 top.pc\[12\] net537 _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ _02652_ _02654_ _02656_ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ _02564_ _02589_ net400 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09212_ _02489_ _02529_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06424_ net812 _01527_ net808 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06355_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__and2_1
X_09143_ _01625_ _04190_ _04193_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout221_A _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _03762_ _03787_ _03814_ _03832_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__or4_1
X_06286_ net1197 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[12\] sky130_fd_sc_hd__and2_1
XFILLER_0_16_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06997__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ top.DUT.register\[1\]\[19\] net703 net643 top.DUT.register\[10\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold720 top.DUT.register\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold731 top.DUT.register\[26\]\[20\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 top.DUT.register\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold753 top.DUT.register\[21\]\[20\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 top.DUT.register\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 top.DUT.register\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06749__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 top.DUT.register\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _01667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 top.DUT.register\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ top.a1.instruction\[7\] top.a1.instruction\[8\] net744 vssd1 vssd1 vccd1
+ vccd1 _04958_ sky130_fd_sc_hd__and3b_1
XANTENNA__07961__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ _02956_ net460 _04008_ net470 _04009_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net279 _02518_ _03355_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_179_Left_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08795__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07809_ net828 _02925_ net468 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o21ai_4
XANTENNA__06921__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ net326 _02090_ _02069_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_28_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ net1398 net260 net494 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10751_ net616 _04977_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__nand2_4
XFILLER_0_55_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13011__RESET_B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ clknet_leaf_32_clk _01016_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net148 net1719 net418 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ clknet_leaf_79_clk top.ru.next_FetchedData\[16\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06762__B _01878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12352_ top.pad.button_control.r_counter\[3\] _06135_ vssd1 vssd1 vccd1 vccd1 _06138_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06988__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ net901 _01382_ _05165_ _05172_ net845 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a311o_1
X_12283_ top.lcd.cnt_20ms\[11\] _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11234_ _05117_ net1242 net402 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10504__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ net925 net1303 net876 _05082_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _04959_ _04965_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nor2_1
X_11096_ net78 _01439_ net848 net1183 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09154__A1 _04169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__B2 _04078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ top.a1.instruction\[10\] net744 top.a1.instruction\[9\] vssd1 vssd1 vccd1
+ vccd1 _04965_ sky130_fd_sc_hd__nand3b_1
XANTENNA__07165__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold80 net101 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold91 _01188_ vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06912__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ clknet_leaf_69_clk _01331_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08992__X _04078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11998_ _05827_ _05828_ _05823_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21oi_1
X_13737_ clknet_leaf_68_clk _00002_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949_ net614 _04986_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13668_ clknet_leaf_90_clk _01209_ net1011 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07401__X _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ clknet_leaf_12_clk _00165_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13599_ clknet_leaf_53_clk _01140_ net1075 vssd1 vssd1 vccd1 vccd1 top.ramload\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08968__B2 _01746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__Q top.a1.instruction\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout507 _04988_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_8
X_09830_ _04825_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10414__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout518 _04983_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_169_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ top.a1.dataIn\[7\] _04765_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_206_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__inv_2
XANTENNA__08886__Y _03977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ _03724_ _03810_ net291 vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__mux2_1
XANTENNA__13682__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _04692_ _04701_ _04694_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07156__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ net397 _02716_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__nor2_1
XANTENNA__13522__RESET_B net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06903__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout171_A _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ net323 net348 _02306_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_25_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ _02641_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1080_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07456_ top.DUT.register\[15\]\[6\] net689 net662 top.DUT.register\[18\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06407_ _01523_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_98_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07387_ top.DUT.register\[26\]\[4\] net722 _02491_ _02503_ vssd1 vssd1 vccd1 vccd1
+ _02504_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _01608_ _01610_ _01723_ _01498_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o22a_1
X_06338_ _01459_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ _03895_ _03916_ _03932_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__and4_1
X_06269_ net1285 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[27\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _03118_ _03120_ _03122_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or4_1
Xhold550 top.DUT.register\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 top.DUT.register\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 top.DUT.register\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 top.DUT.register\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10324__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 top.DUT.register\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12105__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ top.pc\[30\] _04656_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__or2_1
X_12970_ clknet_leaf_118_clk _00516_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11921_ _05734_ _05778_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11852_ _05710_ _05712_ _05709_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09133__B top.a1.instruction\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09439__A2 _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10803_ net191 net1976 net410 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12548__Q top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11783_ _05568_ _05604_ _05632_ _05600_ _05602_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_196_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08111__A2 _03227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ clknet_leaf_105_clk _01068_ net982 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ net206 net2028 net416 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06673__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ clknet_leaf_113_clk _00999_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10665_ net216 net2207 net418 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__mux2_1
X_12404_ clknet_leaf_79_clk top.ru.next_dready net1088 vssd1 vssd1 vccd1 vccd1 top.d_ready
+ sky130_fd_sc_hd__dfrtp_1
X_13384_ clknet_leaf_25_clk _00930_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ net231 net2200 net424 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12335_ _06127_ net743 _06126_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__and3b_1
X_12266_ _06073_ _06085_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11217_ net2322 top.a1.row1\[111\] net405 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__mux2_1
XANTENNA__10234__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__nor2_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11182__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07386__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_208_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11148_ net48 net880 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11079_ net925 _01401_ wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__and3_1
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12458__Q top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_175_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08102__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07310_ _02420_ _02422_ _02424_ _02426_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__or4_4
XFILLER_0_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08290_ _03395_ _03404_ net302 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
XANTENNA__10996__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07241_ top.DUT.register\[18\]\[8\] net778 _02357_ vssd1 vssd1 vccd1 vccd1 _02358_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06664__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10409__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07172_ top.DUT.register\[13\]\[11\] net789 net776 top.DUT.register\[17\]\[11\] _02288_
+ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_200_Left_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09281__A_N _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08810__B1 _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10144__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11173__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07377__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 _01710_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07916__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ _04799_ _04802_ _04810_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net253 net1687 net392 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
X_06956_ top.DUT.register\[10\]\[21\] net727 net776 top.DUT.register\[17\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a22o_1
XANTENNA__07129__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ _04692_ _04694_ _04693_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__o21bai_1
X_06887_ net299 _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout553_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ net476 _02640_ _03728_ net469 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08557_ net281 _03451_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout720_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A _04170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__Y _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ top.DUT.register\[3\]\[14\] net691 net651 top.DUT.register\[17\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
X_08488_ net305 _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07439_ net286 net339 _02428_ _01801_ _02554_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a221o_1
XANTENNA__10319__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ net1682 net150 net512 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__inv_2
X_10381_ net1778 net158 net431 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _05970_ _05977_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__o21a_1
XANTENNA__09409__A _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ top.a1.dataIn\[3\] _05832_ _05881_ top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1
+ _05912_ sky130_fd_sc_hd__or4b_1
XANTENNA__10054__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07368__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 top.DUT.register\[14\]\[16\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net1168 _05021_ net480 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
XANTENNA__07907__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _01511_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_2
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07871__B net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_2
Xfanout893 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_2
X_12953_ clknet_leaf_57_clk _00499_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1080 top.lcd.currentState\[1\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1091 top.DUT.register\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _05690_ _05726_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__nor2_1
X_12884_ clknet_leaf_103_clk _00430_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08883__A3 _03403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11835_ _05694_ _05695_ _05657_ _05687_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06894__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07599__A _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ _05589_ _05623_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__xor2_1
XFILLER_0_184_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13505_ clknet_leaf_45_clk _01051_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net1820 net140 net499 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _05506_ _05557_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13436_ clknet_leaf_17_clk _00982_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10648_ net153 net1810 net375 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09596__A1 _01874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_max_cap351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ clknet_leaf_112_clk _00913_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10579_ net163 top.DUT.register\[19\]\[25\] net504 vssd1 vssd1 vccd1 vccd1 _00723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ top.lcd.cnt_500hz\[7\] _06115_ _06116_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__o21a_1
XANTENNA__07071__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13298_ clknet_leaf_107_clk _00844_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12249_ top.lcd.cnt_20ms\[4\] top.lcd.cnt_20ms\[3\] _06072_ vssd1 vssd1 vccd1 vccd1
+ _06073_ sky130_fd_sc_hd__and3_1
XANTENNA__07359__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire354_A net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10899__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ top.DUT.register\[13\]\[31\] net790 net729 top.DUT.register\[10\]\[31\] _01926_
+ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a221o_1
X_07790_ top.DUT.register\[23\]\[29\] net564 net552 top.DUT.register\[22\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ net307 net301 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__or2_1
X_09460_ _02109_ net840 _04493_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__or3_1
X_06672_ top.DUT.register\[20\]\[1\] net563 net673 top.DUT.register\[19\]\[1\] _01788_
+ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a221o_1
XANTENNA__12475__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07531__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08411_ net1333 net861 net838 _03522_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09391_ _01632_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09808__C1 _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08342_ _03454_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10969__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08273_ _02409_ _02509_ net285 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__mux2_1
XANTENNA__10139__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07224_ top.DUT.register\[25\]\[9\] net713 net709 top.DUT.register\[7\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07155_ top.DUT.register\[9\]\[12\] net716 net752 top.DUT.register\[17\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout301_A _01856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07062__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ net308 net302 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout134 _04230_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout670_A _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 _04923_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout167 net168 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout768_A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _02152_ _03103_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__or2_1
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07770__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ top.a1.dataIn\[0\] net813 _04740_ top.pc\[0\] net457 vssd1 vssd1 vccd1 vccd1
+ _04741_ sky130_fd_sc_hd__a221o_1
X_06939_ top.DUT.register\[14\]\[22\] net793 net751 top.DUT.register\[19\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ net909 top.a1.state\[0\] net908 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or3b_1
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08609_ _02666_ _03712_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_106_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _04614_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11620_ _05470_ _05472_ _05477_ _05479_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11551_ _05393_ _05400_ _05389_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10502_ net209 net1528 net378 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
XANTENNA__09027__B1 _02951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11482_ _05308_ _05330_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ clknet_leaf_47_clk _00767_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10433_ net1635 net219 net509 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ clknet_leaf_12_clk _00698_ net975 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07053__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10364_ net1668 net230 net432 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
X_12103_ _05950_ _05953_ _05955_ _05960_ _05949_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__o41ai_4
XANTENNA__06800__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ clknet_leaf_2_clk _00629_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ net1569 net236 net523 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__mux2_1
X_12034_ _05892_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_148_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10512__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__Y _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _01667_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_4
XANTENNA__07761__B1 _02617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ clknet_leaf_26_clk _00482_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07513__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_8__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12867_ clknet_leaf_34_clk _00413_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11818_ _05647_ net130 vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12798_ clknet_leaf_37_clk _00344_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09805__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _05575_ _05608_ _05574_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07292__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09018__B1 _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ clknet_leaf_4_clk _00965_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_133_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07044__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__C _02611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08960_ net318 _01899_ _01921_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07911_ _03018_ _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__nor2_4
XANTENNA__09336__X _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ _02982_ _03959_ _01982_ _02978_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10422__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ top.DUT.register\[26\]\[26\] net680 net672 top.DUT.register\[19\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07752__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _02883_ _02885_ _02887_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_142_Left_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09512_ _04542_ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_104_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06724_ top.DUT.register\[6\]\[3\] net579 net571 top.DUT.register\[21\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XANTENNA__07016__B _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07504__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _02132_ _04477_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__nand2_1
X_06655_ _01765_ _01767_ _01769_ _01771_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__or4_1
XANTENNA__06858__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09374_ _04412_ _04413_ _04408_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a21oi_1
X_06586_ _01645_ _01653_ _01662_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__and3_1
XFILLER_0_176_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ net296 _03438_ _03401_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_151_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ net464 _03365_ _03371_ _03281_ _03369_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o221a_1
XANTENNA__07283__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07207_ _02309_ _02311_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08187_ net299 _02305_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__nor2_1
XANTENNA__08134__Y _03251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07138_ _02248_ _02250_ _02252_ _02254_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__or4_1
XFILLER_0_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07069_ top.DUT.register\[10\]\[16\] net726 net756 top.DUT.register\[3\]\[16\] _02185_
+ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a221o_1
XANTENNA__11119__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ net146 net1511 net449 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10332__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13770_ clknet_leaf_73_clk _01295_ net1113 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ top.a1.row1\[101\] _04682_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ clknet_leaf_10_clk _00267_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06849__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12652_ clknet_leaf_3_clk _00198_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ _05429_ _05458_ _05432_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__o21a_1
X_12583_ clknet_leaf_52_clk _00129_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11534_ _05389_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__nand2_1
XANTENNA__08471__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07274__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__X _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire332 _02687_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
Xwire343 net344 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
Xwire354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
Xwire365 _02263_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11465_ _05293_ _05295_ _05265_ _05278_ _05285_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_59_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13204_ clknet_leaf_98_clk _00750_ net1005 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07026__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ net1343 net152 net515 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11396_ top.a1.dataIn\[27\] _05255_ _05256_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__and3b_1
XFILLER_0_104_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13135_ clknet_leaf_25_clk _00681_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10347_ net1396 net162 net520 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07982__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ clknet_leaf_116_clk _00612_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08060__X _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ net172 net1842 net435 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__mux2_1
X_12017_ _05873_ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__and2_2
XANTENNA__08526__A2 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12919_ clknet_leaf_111_clk _00465_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06440_ top.a1.instruction\[15\] top.a1.instruction\[16\] net812 _01542_ vssd1 vssd1
+ vccd1 vccd1 _01557_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_192_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06394__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06371_ _01492_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _03217_ _03226_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07787__A _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ _01802_ net272 _03362_ net303 net474 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08041_ _03155_ _03156_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__nand2_2
XANTENNA__06473__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10417__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold902 top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold913 top.DUT.register\[3\]\[26\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07017__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 top.DUT.register\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 top.DUT.register\[16\]\[18\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 top.DUT.register\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 top.DUT.register\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 top.DUT.register\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net218 net1721 net451 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__mux2_1
Xhold979 top.DUT.register\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07973__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ net399 _02928_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10152__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ _03963_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1006_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ top.DUT.register\[13\]\[28\] net676 net648 top.DUT.register\[12\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout466_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ top.DUT.register\[11\]\[31\] net701 net693 top.DUT.register\[3\]\[31\] _02872_
+ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a221o_1
X_06707_ top.DUT.register\[23\]\[4\] net566 net550 top.DUT.register\[4\]\[4\] _01823_
+ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07687_ top.DUT.register\[11\]\[12\] net699 net691 top.DUT.register\[3\]\[12\] _02803_
+ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout633_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09426_ _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__nor2_1
X_06638_ top.DUT.register\[31\]\[2\] net668 net541 top.DUT.register\[5\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09357_ top.pc\[14\] _04368_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06569_ net746 _01647_ _01662_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _03395_ _03400_ _01856_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux2_1
XANTENNA__07256__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09288_ net131 _04322_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09650__B1 _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ _03354_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10327__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11250_ net871 _05112_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and2_1
XANTENNA__07008__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ net210 net1522 net438 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XANTENNA__09953__A1 _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ net367 _01643_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a21oi_1
X_10132_ net210 net1831 net442 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07208__Y _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ net212 net2224 net446 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XANTENNA__10062__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ clknet_leaf_70_clk _01347_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09152__A _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ clknet_leaf_64_clk _01278_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ net1602 net205 net483 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12704_ clknet_leaf_106_clk _00250_ net979 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13684_ clknet_leaf_74_clk net1271 net1089 vssd1 vssd1 vccd1 vccd1 wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ net1997 net218 net406 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ clknet_leaf_0_clk _00181_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ clknet_leaf_76_clk _00112_ net1084 vssd1 vssd1 vccd1 vccd1 top.pc\[31\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07247__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07400__A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06455__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ _05358_ _05376_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10237__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12497_ clknet_leaf_87_clk _00044_ net1082 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08215__B _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 top.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ net327 _05295_ _05273_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_189_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11379_ top.a1.dataIn\[21\] _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__xor2_1
XANTENNA__07955__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ clknet_leaf_38_clk _00664_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13049_ clknet_leaf_55_clk _00595_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07610_ top.DUT.register\[30\]\[11\] net696 net632 top.DUT.register\[27\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10700__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ net463 _03672_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21o_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07541_ top.DUT.register\[23\]\[13\] net564 net659 top.DUT.register\[18\]\[13\] _02657_
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a221o_1
XANTENNA__08132__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ top.a1.instruction\[20\] _01616_ _01640_ top.a1.instruction\[28\] vssd1 vssd1
+ vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08683__B2 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ _02489_ _02529_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__or2_1
X_06423_ top.a1.instruction\[15\] top.a1.instruction\[16\] net812 _01520_ vssd1 vssd1
+ vccd1 vccd1 _01540_ sky130_fd_sc_hd__and4_1
XANTENNA__06694__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ top.a1.instruction\[13\] _01489_ _01716_ _04194_ _01600_ vssd1 vssd1 vccd1
+ vccd1 _04195_ sky130_fd_sc_hd__o311a_1
X_06354_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__and2b_1
XFILLER_0_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07238__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09073_ net310 _03541_ _03843_ _03868_ _03901_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__a2111o_1
X_06285_ net1187 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[11\] sky130_fd_sc_hd__and2_1
XANTENNA__10147__S net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout214_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08024_ _03134_ _03136_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 top.DUT.register\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold721 top.DUT.register\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 top.a1.row2\[10\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09935__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold743 top.DUT.register\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 top.DUT.register\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 top.DUT.register\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 top.DUT.register\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 top.DUT.register\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 top.DUT.register\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ net140 net2105 net393 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout583_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08926_ _04013_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _03058_ net459 _03946_ net470 _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout750_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08795__B _03229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ _02915_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nor2_4
XANTENNA__10610__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ net303 _03534_ _03571_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _02820_ _02284_ _02665_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_0_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ net141 net2026 net417 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07477__A2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09409_ _02175_ _04445_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ net153 net1855 net419 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
XANTENNA__09764__A1_N net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ clknet_leaf_53_clk top.ru.next_FetchedData\[15\] net1078 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12222__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_7__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ top.pad.button_control.r_counter\[3\] _06135_ vssd1 vssd1 vccd1 vccd1 _06137_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10057__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ top.a1.row2\[1\] _05132_ _05166_ _05168_ _05171_ vssd1 vssd1 vccd1 vccd1
+ _05172_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09846__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _06095_ net1117 _06094_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__and3b_1
X_11233_ net871 _05023_ _05036_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ net57 net884 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ net139 net2326 net388 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
X_11095_ net1216 net878 net846 top.ramstore\[13\] vssd1 vssd1 vccd1 vccd1 _01174_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07890__A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ top.a1.instruction\[10\] net744 top.a1.instruction\[9\] vssd1 vssd1 vccd1
+ vccd1 _04964_ sky130_fd_sc_hd__and3b_1
Xhold70 top.DUT.register\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 _01167_ vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 top.a1.row1\[10\] vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
X_13805_ clknet_leaf_69_clk _01330_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11997_ _05850_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13736_ clknet_leaf_69_clk _00001_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__08665__A1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ net2154 net139 net487 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08665__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06676__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_89_clk _01208_ net1013 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10879_ net1585 net150 net490 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ clknet_leaf_118_clk _00164_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ clknet_leaf_53_clk _01139_ net1075 vssd1 vssd1 vccd1 vccd1 top.ramload\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08968__A2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12549_ clknet_leaf_83_clk _00095_ net1007 vssd1 vssd1 vccd1 vccd1 top.pc\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09756__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _01591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07928__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 _04988_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 _04983_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_6
XFILLER_0_158_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _04764_ _04765_ _04198_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__mux2_4
X_06972_ _02079_ _02088_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_206_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _03767_ _03809_ net316 vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__mux2_1
X_09691_ top.edg2.button_i _04705_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__or3_1
XANTENNA__08353__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08642_ _03743_ _03571_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__and2b_1
XANTENNA__09504__B _04525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10430__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ net471 _03675_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08105__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ _02639_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07455_ top.DUT.register\[31\]\[6\] net670 net634 top.DUT.register\[27\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1073_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07311__Y _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ top.a1.instruction\[15\] top.a1.instruction\[16\] _01515_ vssd1 vssd1 vccd1
+ vccd1 _01523_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07386_ top.DUT.register\[14\]\[4\] net794 net586 top.DUT.register\[24\]\[4\] _02502_
+ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a221o_1
XANTENNA__08136__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__inv_2
X_06337_ _01468_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _03837_ _03860_ _03867_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__and4_1
XANTENNA__07092__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06268_ net1456 net895 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[26\] sky130_fd_sc_hd__and2_1
X_08007_ top.DUT.register\[23\]\[21\] net565 net651 top.DUT.register\[17\]\[21\] _03123_
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a221o_1
Xhold540 top.DUT.register\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10605__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06199_ net921 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
Xhold551 top.DUT.register\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 top.DUT.register\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 top.DUT.register\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold584 top.DUT.register\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 top.DUT.register\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12444__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_5_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ top.pc\[30\] _04656_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__nand2_1
X_08909_ net904 top.pc\[27\] _03293_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _02615_ net360 net328 top.a1.dataIn\[23\] net363 vssd1 vssd1 vccd1 vccd1
+ _04880_ sky130_fd_sc_hd__a221o_1
X_11920_ _05739_ _05774_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__xor2_2
XANTENNA__10340__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11851_ _05675_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09133__C top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ net197 net1912 net412 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _05613_ _05641_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_49_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10733_ net211 net1962 net414 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
XANTENNA__13232__RESET_B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__B1 _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ clknet_leaf_7_clk _01067_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_115_clk _00998_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10664_ net221 net2111 net419 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07870__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12403_ clknet_leaf_78_clk net892 net1080 vssd1 vssd1 vccd1 vccd1 top.i_ready sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_52_clk _00929_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10595_ net232 net2124 net424 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12334_ top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] _06123_ vssd1 vssd1 vccd1
+ vccd1 _06127_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09011__A1_N _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06830__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ top.lcd.cnt_20ms\[3\] _06072_ top.lcd.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1
+ _06085_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10515__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11216_ _05039_ _05049_ net369 net404 net1305 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a32o_1
X_12196_ _06035_ _06053_ _06054_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__and3_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__11182__A2 top.pc\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11147_ net922 net1336 net874 _05073_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a31o_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_207_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12874__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output58_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ net26 net863 net835 net1238 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__o22a_1
XANTENNA__10250__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ net203 net1627 net531 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
XANTENNA__07689__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__A1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06897__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08638__B2 _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ clknet_leaf_62_clk _01249_ net1114 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[109\]
+ sky130_fd_sc_hd__dfstp_1
X_07240_ top.DUT.register\[15\]\[8\] net806 net802 top.DUT.register\[31\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a22o_1
XANTENNA__07861__A2 _02977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ top.DUT.register\[28\]\[11\] net739 net585 top.DUT.register\[24\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07074__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08810__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06821__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10425__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout305 _01831_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 _01799_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
X_09812_ _04799_ _04802_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06955_ top.DUT.register\[12\]\[21\] net735 net589 top.DUT.register\[20\]\[21\] _02071_
+ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a221o_1
X_09743_ _03494_ net456 net535 _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout281_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ top.pad.keyCode\[4\] top.pad.keyCode\[6\] top.pad.keyCode\[7\] top.pad.keyCode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_19_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10160__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08877__A1 _03967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06886_ _01993_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_107_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _03532_ _03570_ _03719_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06888__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08556_ net302 _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07507_ top.DUT.register\[24\]\[14\] net544 _02623_ vssd1 vssd1 vccd1 vccd1 _02624_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ _01802_ _03595_ net281 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout713_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07438_ net286 net339 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_102_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07852__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07369_ top.DUT.register\[3\]\[5\] net783 net769 top.DUT.register\[11\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09108_ _02846_ _04160_ _02903_ _02842_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or4b_1
XFILLER_0_150_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07065__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ net1498 net163 net432 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
XANTENNA__07604__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08801__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06812__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09039_ _03283_ net462 _03443_ _03409_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__or4b_1
XANTENNA__10335__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09409__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ _05892_ _05894_ _05884_ _05890_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__a211o_1
Xhold370 top.DUT.register\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 top.DUT.register\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ top.a1.dataIn\[1\] net870 _05019_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_
+ sky130_fd_sc_hd__a22o_1
Xhold392 top.DUT.register\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout850 _05054_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_2
Xfanout861 _01511_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_2
Xfanout872 _04677_ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout883 _01439_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10070__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ clknet_leaf_33_clk _00498_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1070 top.DUT.register\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 top.DUT.register\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net125 net126 _05747_ _05755_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a211o_1
XANTENNA__06879__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1092 top.DUT.register\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_12883_ clknet_leaf_109_clk _00429_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11834_ top.a1.dataIn\[7\] _05625_ _05654_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__or3b_1
XFILLER_0_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11765_ top.a1.dataIn\[8\] _05623_ _05624_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08096__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10716_ top.DUT.register\[23\]\[30\] net144 net499 vssd1 vssd1 vccd1 vccd1 _00856_
+ sky130_fd_sc_hd__mux2_1
X_13504_ clknet_leaf_13_clk _01050_ net968 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ _05483_ _05505_ _05486_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07843__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13435_ clknet_leaf_2_clk _00981_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10647_ net157 net1734 net375 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ clknet_leaf_104_clk _00912_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09596__A2 _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ net166 net2168 net503 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__mux2_1
XANTENNA__08063__X _03180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ top.lcd.cnt_500hz\[7\] _06115_ net743 vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__a21boi_1
X_13297_ clknet_leaf_9_clk _00843_ net971 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_197_Left_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08998__X _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ top.lcd.cnt_20ms\[2\] top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] vssd1 vssd1
+ vccd1 vccd1 _06072_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ _06023_ _06026_ _06028_ _06039_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__o31a_1
XANTENNA__08020__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__A0 _03395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__Y _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ net307 net301 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08859__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06671_ top.DUT.register\[22\]\[1\] net554 net657 top.DUT.register\[28\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ net904 top.pc\[5\] _03291_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a22o_1
X_09390_ _04426_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08341_ _02849_ _03453_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07295__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08272_ _02367_ _02470_ net313 vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07223_ _02334_ _02336_ _02338_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__or4_2
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07047__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07154_ top.DUT.register\[22\]\[12\] net604 net756 top.DUT.register\[3\]\[12\] _02270_
+ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a221o_1
XANTENNA__07598__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07085_ net305 net282 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__nor2_1
XANTENNA__10155__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08701__X _03801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout496_A _04999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout135 _04208_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_4
Xfanout146 _04950_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _04923_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_1
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_2
X_07987_ _02152_ _03103_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__and2_1
Xfanout179 _04867_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__Y _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ top.DUT.register\[21\]\[22\] net609 net601 top.DUT.register\[5\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a22o_1
X_09726_ _04199_ _04735_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__and2_1
X_09657_ net909 top.a1.state\[0\] net908 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__nor3b_1
X_06869_ top.DUT.register\[8\]\[25\] net594 net769 top.DUT.register\[11\]\[25\] _01985_
+ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08608_ _02821_ _03691_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2b_1
X_09588_ top.pc\[27\] _04583_ top.pc\[28\] vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08539_ _03627_ _03643_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_46_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08078__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07987__X _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _05389_ net248 vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__and2_1
XANTENNA__07825__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10501_ net213 net1788 net378 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ top.a1.dataIn\[16\] _05338_ _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05342_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09027__B2 _04082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ clknet_leaf_31_clk _00766_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10432_ net1525 net227 net509 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13151_ clknet_leaf_32_clk _00697_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10363_ net1403 net233 net432 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
X_12102_ _05950_ _05953_ _05955_ _05960_ _05949_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__o41a_2
X_13082_ clknet_leaf_16_clk _00628_ net987 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08611__X _03715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ net1381 net245 net523 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__mux2_1
X_12033_ _05860_ _05863_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08002__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09750__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07761__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__A2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _01675_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
Xfanout691 net694 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ clknet_leaf_44_clk _00481_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12866_ clknet_leaf_11_clk _00412_ net976 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11817_ _05640_ net130 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_56_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12797_ clknet_leaf_0_clk _00343_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08218__B _02132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07277__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ _05575_ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07816__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__RESET_B net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10820__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09018__B2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _05536_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07029__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13418_ clknet_leaf_118_clk _00964_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ clknet_leaf_39_clk _00895_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07910_ _03020_ _03022_ _03024_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__or4_1
XANTENNA__10703__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ net1268 net861 net838 _03980_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__a22o_1
XANTENNA__07201__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ _02906_ _02932_ _02956_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__or3_1
X_07772_ top.DUT.register\[23\]\[30\] net566 net654 top.DUT.register\[17\]\[30\] _02888_
+ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a221o_1
X_06723_ top.DUT.register\[5\]\[3\] net543 net642 top.DUT.register\[9\]\[3\] _01839_
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a221o_1
X_09511_ _02047_ _02616_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11836__B1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12592__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _02132_ _04477_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06654_ top.DUT.register\[21\]\[2\] net569 net549 top.DUT.register\[4\]\[2\] _01770_
+ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ _02222_ _04411_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09257__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06585_ net747 _01656_ _01658_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__and3_1
XANTENNA__09257__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ _03345_ _03351_ _01800_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__B2 top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ _01736_ _03288_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__or2_4
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout411_A _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A _04987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ top.DUT.register\[27\]\[10\] net770 _02307_ _02322_ vssd1 vssd1 vccd1 vccd1
+ _02323_ sky130_fd_sc_hd__a211o_1
X_08186_ _03298_ _03301_ net320 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07137_ top.DUT.register\[21\]\[13\] net608 net715 top.DUT.register\[9\]\[13\] _02253_
+ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07068_ top.DUT.register\[25\]\[16\] net711 net707 top.DUT.register\[7\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10613__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06599__A top.a1.instruction\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _01409_ _01643_ net138 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a21oi_1
X_10981_ net1486 net141 net483 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ clknet_leaf_116_clk _00266_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12651_ clknet_leaf_3_clk _00197_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_0__f_clk_X clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07259__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11055__A1 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ _05459_ _05462_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_176_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ clknet_leaf_48_clk _00128_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11533_ _05392_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_4
Xwire355 _01961_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11464_ _05280_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire366 net368 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13203_ clknet_leaf_107_clk _00749_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10415_ net1588 net156 net513 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__A0 _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ top.a1.dataIn\[26\] _05250_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ net1374 net168 net520 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13134_ clknet_leaf_94_clk _00680_ net999 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06785__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_27_clk _00611_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ net176 net1612 net435 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__mux2_1
XANTENNA__10523__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _05830_ _05864_ _05844_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_206_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07734__A1 _02612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ clknet_leaf_103_clk _00464_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_192_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12849_ clknet_leaf_10_clk _00395_ net972 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06370_ net34 top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__nand2_1
XANTENNA__08516__X _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_211_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 top.DUT.register\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold914 top.DUT.register\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 top.DUT.register\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 top.a1.row1\[108\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 top.DUT.register\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 top.DUT.register\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13516__RESET_B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold969 top.DUT.register\[8\]\[23\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net221 net1840 net451 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__mux2_1
XANTENNA__06776__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11__f_clk_X clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _02203_ _03871_ _04029_ net274 _04026_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o221a_1
XANTENNA__10433__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08873_ _02983_ _03962_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout194_A _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07824_ _02934_ _02936_ _02938_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__or4_1
XFILLER_0_169_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07755_ top.DUT.register\[30\]\[31\] net697 net629 top.DUT.register\[29\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout361_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06866__B _01981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout459_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ top.DUT.register\[22\]\[4\] net554 net543 top.DUT.register\[5\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a22o_1
X_07686_ top.DUT.register\[15\]\[12\] net687 net667 top.DUT.register\[31\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09425_ _04443_ _04447_ _04446_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__o21ai_2
X_06637_ net826 _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__or2_2
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__B2 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06568_ top.DUT.register\[19\]\[0\] net672 net668 top.DUT.register\[31\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__a22o_1
X_09356_ _04394_ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07330__X _02447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ _03420_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ net135 _04328_ _04331_ net821 net915 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10608__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06499_ _01595_ net854 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__nand2_2
XFILLER_0_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08238_ net296 _03353_ _03349_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o21a_1
XANTENNA__07661__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08169_ _02827_ _03060_ _03259_ _03285_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__or4_2
XFILLER_0_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ net214 net1696 net438 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07413__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ _01386_ net822 _04210_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10131_ net213 net1752 net442 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__mux2_1
XANTENNA__10343__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10062_ net216 net1786 net446 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07192__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ clknet_leaf_70_clk _01346_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13752_ clknet_leaf_64_clk _01277_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ net1469 net209 net482 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XANTENNA__12821__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06495__C top.a1.instruction\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12703_ clknet_leaf_23_clk _00249_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ clknet_leaf_75_clk _01224_ net1091 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10895_ net1577 net220 net407 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07888__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12225__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ clknet_leaf_19_clk _00180_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10518__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ clknet_leaf_76_clk _00111_ net1084 vssd1 vssd1 vccd1 vccd1 top.pc\[30\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_156_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11516_ _05358_ _05376_ _05361_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12496_ clknet_leaf_88_clk _00043_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ _05306_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ _05228_ _05230_ top.a1.dataIn\[20\] vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06758__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10329_ net1508 net238 net519 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__mux2_1
X_13117_ clknet_leaf_118_clk _00663_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13048_ clknet_leaf_33_clk _00594_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07183__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07540_ top.DUT.register\[10\]\[13\] net643 net623 top.DUT.register\[16\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07471_ _02489_ _02549_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06973__Y _02090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09210_ _01808_ net337 _04249_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o21a_1
X_06422_ net809 _01518_ _01536_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__and3_1
XANTENNA__12216__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net912 _01597_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__xnor2_1
X_06353_ top.pad.count\[1\] top.pad.count\[0\] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__and2b_1
XFILLER_0_174_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10428__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13768__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ _03589_ _03608_ _03656_ _03631_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__or4b_1
X_06284_ net2232 net899 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[10\] sky130_fd_sc_hd__and2_1
XANTENNA__07643__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08023_ top.DUT.register\[21\]\[19\] net568 _03137_ _03139_ vssd1 vssd1 vccd1 vccd1
+ _03140_ sky130_fd_sc_hd__a211o_1
XANTENNA__06997__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold700 top.DUT.register\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold711 top.DUT.register\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 top.DUT.register\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold733 top.DUT.register\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 top.DUT.register\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09518__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 top.DUT.register\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold766 top.DUT.register\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06749__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold777 top.DUT.register\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold788 top.DUT.register\[24\]\[28\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 top.DUT.register\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _04079_ _04737_ net536 _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout1116_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _02957_ _04012_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout576_A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _03928_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nand2_1
XANTENNA__07174__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__A _02366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _02917_ _02919_ _02921_ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or4_1
X_08787_ _03232_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06921__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _02743_ _02853_ _02854_ _02823_ _02666_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_0_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout910_A net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07669_ top.DUT.register\[30\]\[10\] net695 net655 top.DUT.register\[28\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _02175_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12207__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ net154 net1755 net418 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07501__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ _04379_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__nand2_1
XANTENNA__10338__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ _06135_ _06136_ net814 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__and3b_1
XANTENNA__07634__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06988__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ top.a1.row2\[25\] _05134_ _05138_ top.a1.row2\[9\] _05170_ vssd1 vssd1 vccd1
+ vccd1 _05171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12281_ top.lcd.cnt_20ms\[10\] top.lcd.cnt_20ms\[9\] _06091_ vssd1 vssd1 vccd1 vccd1
+ _06095_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _05116_ net1484 net402 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ net925 net1351 net876 _05081_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a31o_1
X_10114_ net143 net1963 net389 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ net76 net879 net847 net1184 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
X_10045_ net139 net1783 net531 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XANTENNA__10801__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 _01171_ vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 top.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 top.ramload\[4\] vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net86 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12301__B _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ clknet_leaf_69_clk _01329_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _05851_ _05852_ _05854_ _05855_ _05805_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_67_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13735_ clknet_leaf_69_clk _00000_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10947_ net1419 net143 net488 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09862__A1 _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07873__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_90_clk _01207_ net1012 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
X_10878_ net1378 net156 net490 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12617_ clknet_leaf_27_clk _00163_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10248__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ clknet_leaf_56_clk _01138_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramload\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12548_ clknet_leaf_83_clk _00094_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06979__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ clknet_leaf_89_clk _00026_ net1015 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09338__A _02264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06314__X _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout509 _04987_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _02083_ _02084_ _02085_ _02087_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_206_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _02154_ _02176_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__or2_1
XANTENNA__10711__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ _04691_ _04699_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nor2_1
XANTENNA__07156__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1080 net1081 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
X_08641_ net274 _03552_ _03556_ net269 vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__a2bb2o_1
Xfanout1091 net1121 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06903__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08572_ net477 _02821_ _02823_ net458 _03676_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07523_ _02243_ _02638_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_25_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout157_A _04923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07454_ top.DUT.register\[1\]\[6\] net705 net563 top.DUT.register\[20\]\[6\] _02570_
+ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09520__B _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06405_ net809 _01521_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__nor2_1
XANTENNA__10158__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07385_ top.DUT.register\[23\]\[4\] net732 net751 top.DUT.register\[19\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06419__A1 top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06336_ _01331_ _01330_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07616__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ _01618_ _04174_ _04175_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__or4_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09055_ _03779_ _03798_ _03808_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__and4_1
X_06267_ net1324 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[25\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ top.DUT.register\[6\]\[21\] net577 net624 top.DUT.register\[16\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a22o_1
Xhold530 top.DUT.register\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09908__A2 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06198_ net36 net35 net38 net37 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nor4_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08152__A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold541 top.DUT.register\[29\]\[2\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold552 top.DUT.register\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 top.DUT.register\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12526__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 top.DUT.register\[24\]\[17\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 top.DUT.register\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold596 top.DUT.register\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__B2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ net149 net1968 net390 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _03996_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nor2_1
XANTENNA__10621__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ net819 _04534_ _04535_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__or3_1
XANTENNA__08344__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ _03930_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12413__RESET_B net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__A top.a1.instruction\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _05631_ _05635_ net130 _05637_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09133__D top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10801_ net200 net2118 net410 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11781_ _05613_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__or2_1
XANTENNA__09844__A1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11100__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13520_ clknet_leaf_117_clk _01066_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06658__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ net214 net1841 net414 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
XANTENNA__07855__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13619__RESET_B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13451_ clknet_leaf_6_clk _00997_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10663_ net224 top.DUT.register\[22\]\[10\] net418 vssd1 vssd1 vccd1 vccd1 _00804_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10068__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12402_ clknet_leaf_60_clk top.a1.nextHex\[7\] net1102 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09857__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ net238 net1705 net424 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__mux2_1
X_13382_ clknet_leaf_49_clk _00928_ net1048 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12333_ top.lcd.cnt_500hz\[12\] _06123_ top.lcd.cnt_500hz\[13\] vssd1 vssd1 vccd1
+ vccd1 _06126_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_12264_ _06080_ _06084_ net1117 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_186_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11215_ _05035_ _05046_ _05108_ net404 net1186 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a32o_1
XANTENNA__08032__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ _06053_ _06054_ _06035_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a21oi_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__08997__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07386__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
XANTENNA__08583__B2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__B1 _04359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
X_11146_ net47 net880 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_207_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10531__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__B _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11077_ net25 net852 _05054_ net1524 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10028_ net209 net1386 net530 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
XANTENNA__07406__A _02517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_201_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11979_ _05813_ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__xnor2_1
X_13718_ clknet_leaf_62_clk _01248_ net1109 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07846__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ clknet_leaf_110_clk net1226 net995 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09767__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07170_ top.DUT.register\[29\]\[11\] net785 net731 top.DUT.register\[23\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_120_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10706__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
XANTENNA__08574__A1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07377__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
X_09811_ _04808_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand2_1
XANTENNA__11173__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
XANTENNA__10441__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ top.pc\[4\] net817 net457 _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_1
X_06954_ top.DUT.register\[28\]\[21\] net739 net793 top.DUT.register\[14\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07129__A2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09673_ _04691_ _04692_ _01480_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_207_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06885_ _01995_ _01997_ _01999_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__or4_4
X_08624_ net306 _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08555_ _03562_ _03660_ net295 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout441_A _04976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09287__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout539_A _03291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07506_ top.DUT.register\[26\]\[14\] net679 net639 top.DUT.register\[9\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_194_Right_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08486_ _03484_ _03594_ net289 vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07437_ _02553_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ top.DUT.register\[13\]\[5\] net791 net595 top.DUT.register\[8\]\[5\] _02484_
+ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09107_ net475 _04159_ _02880_ _03417_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__or4b_1
XFILLER_0_134_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06319_ top.lcd.nextState\[0\] top.lcd.currentState\[0\] _01453_ vssd1 vssd1 vccd1
+ vccd1 _01458_ sky130_fd_sc_hd__mux2_1
X_07299_ top.DUT.register\[1\]\[1\] net780 net763 top.DUT.register\[30\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a22o_1
XANTENNA__10616__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_135_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09038_ _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 top.DUT.register\[7\]\[7\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 top.DUT.register\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07368__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 top.DUT.register\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ top.a1.halfData\[1\] _05008_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or2_1
Xhold393 top.DUT.register\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__B2 _03670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _02613_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_8
Xfanout851 _05052_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_2
Xfanout862 _05053_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_2
XANTENNA__10351__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 _04224_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout895 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_2
X_12951_ clknet_leaf_112_clk _00497_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1060 top.DUT.register\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1071 top.DUT.register\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net125 net126 _05728_ _05747_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a211o_1
Xhold1082 top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 top.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_104_clk _00428_ net983 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09441__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11833_ _05682_ _05686_ _05658_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_64_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09160__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ _05623_ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13503_ clknet_leaf_23_clk _01049_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10715_ net1999 net148 net497 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11695_ _05535_ _05541_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13434_ clknet_leaf_15_clk _00980_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ net160 net1582 net376 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10526__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__B1 _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ clknet_leaf_82_clk _00911_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10577_ net172 net2167 net502 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _06115_ net742 _06114_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ clknet_leaf_115_clk _00842_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08005__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ net1149 _05994_ net612 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07359__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__B1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12178_ _06023_ _06026_ _06031_ _06028_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08520__A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07407__Y _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net924 net1293 net876 _05064_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a31o_1
XANTENNA__10261__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06319__A0 top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ _01780_ _01782_ _01784_ _01786_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__or4_1
XANTENNA__07531__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A _02244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08340_ _02849_ _03453_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07819__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08271_ _03384_ _03385_ net291 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ top.DUT.register\[22\]\[9\] net606 net731 top.DUT.register\[23\]\[9\] _02328_
+ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__a221o_1
X_07153_ top.DUT.register\[14\]\[12\] net792 net754 top.DUT.register\[18\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkload59_A clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10436__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A2 _02714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _02028_ _02200_ net282 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1029_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout125 _05758_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
XANTENNA_fanout391_A _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _04208_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
Xfanout147 _04941_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout489_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 _04913_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout169 _04895_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
X_07986_ net825 _03102_ _02617_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07770__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ top.a1.instruction\[11\] _04729_ _04738_ net34 net745 vssd1 vssd1 vccd1 vccd1
+ _04739_ sky130_fd_sc_hd__o311a_2
X_06937_ top.DUT.register\[17\]\[22\] net776 _02053_ vssd1 vssd1 vccd1 vccd1 _02054_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout656_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ net908 net909 top.a1.state\[0\] _04676_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__and4b_1
XFILLER_0_179_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06868_ top.DUT.register\[10\]\[25\] net728 net772 top.DUT.register\[27\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08607_ net397 _02663_ _03706_ net472 _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__o221a_1
XANTENNA__09010__A1_N _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ top.pc\[27\] top.pc\[28\] _04583_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06799_ top.DUT.register\[21\]\[30\] net610 net722 top.DUT.register\[26\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA__06730__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12714__CLK clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08538_ _02522_ _03630_ _03642_ net464 _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_46_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _03577_ _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ net218 net1771 net378 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
XANTENNA__09025__A1_N _02977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09027__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__and2_1
XFILLER_0_190_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ net1815 net230 net511 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XANTENNA__10346__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07589__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ clknet_leaf_38_clk _00696_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ net2085 net236 net432 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XANTENNA__06797__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12101_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10293_ net2004 net250 net524 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__mux2_1
X_13081_ clknet_leaf_56_clk _00627_ net1094 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08538__A1 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _05861_ _05862_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__and2_1
XANTENNA__09735__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 _01185_ vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06412__X _01529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _01684_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_2
XANTENNA__07761__A2 _02877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__X _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 _01675_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout692 net694 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_4
XANTENNA__09499__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__B _04078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ clknet_leaf_22_clk _00480_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13634__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07513__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12865_ clknet_leaf_45_clk _00411_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06721__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11816_ _05639_ _05605_ _05675_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12796_ clknet_leaf_18_clk _00342_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11747_ _05571_ _05580_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _05520_ _05529_ _05533_ _05525_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13417_ clknet_leaf_28_clk _00963_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10256__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ net229 net2094 net376 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XANTENNA__12037__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09974__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13348_ clknet_leaf_29_clk _00894_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06788__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__Y _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13279_ clknet_leaf_22_clk _00825_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_47_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08250__A _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07840_ _02956_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07752__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ top.DUT.register\[1\]\[30\] net706 net571 top.DUT.register\[21\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06960__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _02047_ _02616_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_1
X_06722_ top.DUT.register\[11\]\[3\] net702 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07504__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08701__B2 _03800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ net840 _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__nor2_2
X_06653_ top.DUT.register\[3\]\[2\] net692 net688 top.DUT.register\[15\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_56_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ _02222_ _04411_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06584_ net747 _01653_ _01658_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__and3_4
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08323_ _01856_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_A _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08254_ _01736_ _03288_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07205_ top.DUT.register\[6\]\[10\] net596 net750 top.DUT.register\[19\]\[10\] _02321_
+ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1087_A top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ _03299_ _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07136_ top.DUT.register\[13\]\[13\] net788 net719 top.DUT.register\[26\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06779__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07067_ top.DUT.register\[28\]\[16\] net738 net734 top.DUT.register\[12\]\[16\] _02183_
+ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a221o_1
XANTENNA__11119__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ top.DUT.register\[8\]\[18\] net556 net659 top.DUT.register\[18\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__Y _02003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _04210_ _04211_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o21a_1
X_10980_ net1543 net143 net484 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XANTENNA__08159__X _03276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09639_ _04209_ _04221_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13045__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12650_ clknet_leaf_116_clk _00196_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ _05420_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ clknet_leaf_39_clk _00127_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11532_ _05345_ _05381_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire345 _02389_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10076__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _05248_ _05255_ net478 _05256_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_83_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ clknet_leaf_107_clk _00748_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09956__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ top.DUT.register\[14\]\[26\] net158 net514 vssd1 vssd1 vccd1 vccd1 _00564_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11394_ _05225_ _05232_ _05233_ _01393_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a22o_2
XFILLER_0_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ clknet_leaf_113_clk _00679_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10345_ net1757 net171 net517 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XANTENNA__10804__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07982__A2 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ clknet_leaf_24_clk _00610_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10276_ net180 net1730 net435 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__mux2_1
XANTENNA__12304__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ _05873_ _05875_ _05868_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07195__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06942__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12917_ clknet_leaf_101_clk _00463_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12848_ clknet_leaf_116_clk _00394_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12779_ clknet_leaf_4_clk _00325_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06473__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09775__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold904 top.DUT.register\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 top.DUT.register\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 top.a1.hexop\[2\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold937 top.DUT.register\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold948 top.pad.keyCode\[1\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 top.DUT.register\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ net223 top.DUT.register\[2\]\[10\] net450 vssd1 vssd1 vccd1 vccd1 _00164_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10714__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _03942_ _04028_ net293 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08872_ _02983_ _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_209_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13556__RESET_B net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07186__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07823_ top.DUT.register\[11\]\[28\] net701 net565 top.DUT.register\[23\]\[28\] _02939_
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06933__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout187_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ top.DUT.register\[22\]\[31\] net554 net547 top.DUT.register\[24\]\[31\] _02870_
+ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06705_ top.DUT.register\[15\]\[4\] net689 net669 top.DUT.register\[31\]\[4\] _01821_
+ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07685_ top.DUT.register\[7\]\[12\] net572 net568 top.DUT.register\[21\]\[12\] _02801_
+ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1096_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09424_ _02152_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__xor2_1
X_06636_ net855 _01752_ _01751_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12234__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ _04380_ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and2_1
XANTENNA__08438__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06567_ _01645_ _01656_ _01662_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__and3_2
XFILLER_0_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ net475 _02842_ net462 _03409_ _03415_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__o221a_1
XANTENNA__08989__A1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09286_ _04329_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07110__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06498_ net841 net856 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08237_ net319 _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ _02845_ _02849_ _03283_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07119_ top.DUT.register\[19\]\[14\] net765 net708 top.DUT.register\[7\]\[14\] _02235_
+ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a221o_1
XANTENNA__09261__A_N _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ top.DUT.register\[20\]\[22\] net561 _03213_ _03215_ vssd1 vssd1 vccd1 vccd1
+ _03216_ sky130_fd_sc_hd__a211o_1
X_10130_ net216 net2059 net442 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ net221 net1615 net447 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
XANTENNA__07177__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06924__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_70_clk _01345_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ clknet_leaf_65_clk _01276_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10963_ net1866 net214 net481 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_82_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12702_ clknet_leaf_38_clk _00248_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09720__Y _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13682_ clknet_leaf_75_clk _01223_ net1090 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
X_10894_ net1998 net226 net406 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12633_ clknet_leaf_61_clk _00179_ net1101 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08429__B1 _03371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ clknet_leaf_87_clk _00110_ net1018 vssd1 vssd1 vccd1 vccd1 top.pc\[29\] sky130_fd_sc_hd__dfstp_1
XANTENNA__08065__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13679__Q net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07101__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A2 _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11515_ _05352_ _05354_ _05363_ _05364_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_156_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06455__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ clknet_leaf_90_clk _00042_ net1011 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11446_ _05269_ _05303_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10534__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11377_ _05235_ _05237_ top.a1.dataIn\[22\] _05231_ vssd1 vssd1 vccd1 vccd1 _05238_
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_21_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07955__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13116_ clknet_leaf_101_clk _00662_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ net1352 net244 net519 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__mux2_1
X_13047_ clknet_leaf_107_clk _00593_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ net253 net2150 net436 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__X _01717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08132__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ _02567_ _02586_ net826 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_2
XFILLER_0_158_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07340__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06421_ net811 _01521_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06694__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09140_ net912 _01513_ _01601_ _01632_ net817 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__a311o_1
X_06352_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__nor2_1
XFILLER_0_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06283_ net1653 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[9\] sky130_fd_sc_hd__and2_1
X_09071_ _03675_ _03700_ _03728_ _03748_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_20_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08022_ top.DUT.register\[2\]\[19\] net683 net548 top.DUT.register\[4\]\[19\] _03138_
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 top.DUT.register\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top.DUT.register\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold723 top.DUT.register\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 top.DUT.register\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10444__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold745 top.DUT.register\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 top.DUT.register\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 top.DUT.register\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 top.DUT.register\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _04171_ _04662_ _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_139_Left_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold789 top.DUT.register\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ _02957_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__or2_1
XANTENNA__07159__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ net477 _03055_ _03054_ net399 vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout569_A _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07806_ top.DUT.register\[20\]\[29\] net560 net623 top.DUT.register\[16\]\[29\] _02922_
+ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09253__B _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ _03130_ _03864_ _03131_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07737_ _02796_ _02326_ _02744_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_0_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08123__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07668_ _02778_ _02780_ _02782_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_148_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ net857 _02525_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__a21oi_4
X_06619_ _01719_ _01735_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__nand2_4
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ _02223_ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ _02264_ _04378_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__nand2_1
XANTENNA__07501__B _02615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _04313_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ top.a1.row1\[57\] _05140_ _05149_ top.a1.row1\[105\] _05169_ vssd1 vssd1
+ vccd1 vccd1 _05170_ sky130_fd_sc_hd__a221o_1
X_12280_ top.lcd.cnt_20ms\[9\] top.lcd.cnt_20ms\[8\] _06090_ top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11231_ net871 _05018_ _05033_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ net56 net884 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__and2_1
X_10113_ net148 net2304 net386 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ net75 net878 net846 net1194 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a22o_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net145 net2078 net531 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XANTENNA__06420__X _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 _01187_ vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 net104 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 net83 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net113 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _01182_ vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09731__X _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ clknet_leaf_69_clk _01328_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11995_ _05854_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_55_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13734_ clknet_leaf_62_clk _01264_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_10946_ net1966 net148 net485 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07322__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06676__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13665_ clknet_leaf_90_clk _01206_ net1010 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
X_10877_ net1481 net159 net490 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
XANTENNA__10529__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ clknet_leaf_25_clk _00162_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13596_ clknet_leaf_55_clk _01137_ net1095 vssd1 vssd1 vccd1 vccd1 top.ramload\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11957__B1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12547_ clknet_leaf_83_clk _00093_ net1009 vssd1 vssd1 vccd1 vccd1 top.pc\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12478_ clknet_leaf_89_clk _00025_ net1015 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09378__B2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10264__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ _05248_ _05257_ net478 _05254_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09338__B _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07389__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ top.DUT.register\[5\]\[21\] net601 net593 top.DUT.register\[8\]\[21\] _02086_
+ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1070 net1072 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_4
X_08640_ net462 _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_1
Xfanout1081 net1091 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12478__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ net397 _02822_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08105__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07522_ _02243_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07313__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07602__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload89_A clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ top.DUT.register\[7\]\[6\] net575 net698 top.DUT.register\[30\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XANTENNA__10439__S net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06404_ _01518_ _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07384_ _02494_ _02496_ _02498_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__or4_1
X_09123_ top.a1.instruction\[12\] _01603_ _01608_ vssd1 vssd1 vccd1 vccd1 _04176_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_98_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06335_ net1118 _01458_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1059_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ _03713_ _03736_ _03756_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07092__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06266_ top.ramload\[24\] net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08005_ top.DUT.register\[14\]\[21\] net664 net656 top.DUT.register\[28\]\[21\] _03121_
+ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold520 top.DUT.register\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10174__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06197_ net2075 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold531 top.DUT.register\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 top.DUT.register\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold553 top.DUT.register\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 top.DUT.register\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 top.DUT.register\[30\]\[7\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 top.DUT.register\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _01670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 top.DUT.register\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10902__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _04039_ net455 net534 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__o211a_4
XTAP_TAPCELL_ROW_51_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ _03995_ _03978_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__and2b_1
X_09887_ net174 net1882 net391 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08838_ _03032_ _03180_ _03914_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08769_ _03132_ _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10800_ net203 net2045 net412 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__mux2_1
X_11780_ _05594_ _05596_ _05606_ _05615_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07304__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11100__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ net217 net1290 net414 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
XANTENNA__10349__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__A2 _01773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ clknet_leaf_118_clk _00996_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ net228 net1814 net420 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ clknet_leaf_60_clk _00009_ net1102 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13381_ clknet_leaf_39_clk _00927_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ net246 net1703 net425 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ top.lcd.cnt_500hz\[12\] _06123_ _06125_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__o21a_1
X_12263_ top.lcd.cnt_20ms\[3\] _06072_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__xor2_1
XANTENNA__10084__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09158__B _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08062__B _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11214_ _05032_ _05044_ _05108_ net404 net1248 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_186_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12194_ _06053_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__nand2_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__09780__A1 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
X_11145_ net923 net1327 net875 _05072_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10812__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07791__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_207_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net23 net863 net835 net1196 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__o22a_1
X_10027_ net215 net2340 net529 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
XANTENNA__07406__B _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06897__A2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_201_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _05811_ _05821_ _05833_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13717_ clknet_leaf_65_clk _01247_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10929_ net1785 net217 net485 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__mux2_1
XANTENNA__06649__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__S net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_88_clk net1314 net1016 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09599__A1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13579_ clknet_leaf_63_clk _01120_ net1107 vssd1 vssd1 vccd1 vccd1 top.a1.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10602__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07074__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06821__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08540__X _03647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout307 _01831_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
X_09810_ _01414_ _04411_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__nand2_1
XANTENNA__08574__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10722__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout318 net319 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 _04820_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
X_09741_ net820 _04241_ top.a1.dataIn\[4\] net813 vssd1 vssd1 vccd1 vccd1 _04751_
+ sky130_fd_sc_hd__a2bb2o_1
X_06953_ _02049_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08326__A2 _03439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ top.pad.keyCode\[1\] top.pad.keyCode\[0\] top.pad.keyCode\[2\] top.pad.keyCode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__or4b_2
X_06884_ top.DUT.register\[13\]\[25\] net791 net779 top.DUT.register\[18\]\[25\] _02000_
+ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a221o_1
XANTENNA__07534__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__X _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ _03538_ _03725_ net282 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__mux2_1
XANTENNA__06888__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout267_A _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08554_ net320 _03610_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o21ai_1
X_07505_ top.DUT.register\[14\]\[14\] net663 net635 top.DUT.register\[25\]\[14\] _02621_
+ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a221o_1
XANTENNA__07332__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ _03536_ _03593_ net313 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__mux2_1
XANTENNA__10169__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A0 top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ _01738_ net285 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07367_ top.DUT.register\[5\]\[5\] net602 net590 top.DUT.register\[20\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout601_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _02830_ _02836_ _03180_ _03229_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__or4b_1
XFILLER_0_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06318_ _01448_ _01454_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07065__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07298_ top.DUT.register\[6\]\[1\] net598 net714 top.DUT.register\[25\]\[1\] _02414_
+ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _04085_ _04088_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__nand2_1
XANTENNA__06812__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06249_ top.ramload\[7\] net893 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[7\]
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_211_Right_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold350 top.DUT.register\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 top.DUT.register\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 top.DUT.register\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 top.DUT.register\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10632__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 top.DUT.register\[4\]\[26\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09706__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 _01515_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_2
Xfanout841 _01594_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
Xfanout852 _05052_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_1
X_09939_ net818 _04616_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06411__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 _05053_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout874 net876 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_2
X_12950_ clknet_leaf_102_clk _00496_ net984 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09514__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_2
Xhold1050 top.DUT.register\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net125 net126 _05747_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a21oi_2
Xhold1061 top.DUT.register\[20\]\[9\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__B top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1072 top.DUT.register\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 top.pad.keyCode\[5\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06879__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12881_ clknet_leaf_7_clk _00427_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1094 top.DUT.register\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_11832_ _05663_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_64_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11763_ top.a1.dataIn\[9\] _05612_ _05614_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__and3_1
XANTENNA__10079__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13502_ clknet_leaf_38_clk _01048_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10714_ net1407 net152 net500 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
X_11694_ _05549_ _05551_ _05553_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ clknet_leaf_43_clk _00979_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ net164 net1953 net377 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
XANTENNA__10807__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13493__RESET_B net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13364_ clknet_leaf_96_clk _00910_ net1002 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08253__B2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10576_ net176 net1960 net502 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__mux2_1
X_12315_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] top.lcd.cnt_500hz\[6\] _01447_
+ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ clknet_leaf_20_clk _00841_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06305__B net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ _06006_ net612 _06071_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06555__C_N top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12177_ _06026_ _06031_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__or2_1
XANTENNA__10542__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11128_ net69 net882 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11059_ net5 net862 net834 net1197 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__o22a_1
XANTENNA__11312__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09632__A _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09351__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08248__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09808__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ _02285_ _02327_ net313 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__mux2_1
XANTENNA__07295__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10784__Y _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07221_ top.DUT.register\[5\]\[9\] net602 net728 top.DUT.register\[10\]\[9\] _02337_
+ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a221o_1
XANTENNA__10717__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07152_ top.DUT.register\[23\]\[12\] net730 net759 top.DUT.register\[2\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a22o_1
XANTENNA__07047__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07083_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10452__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout126 _05759_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07755__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _04208_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
X_07985_ _03088_ _03092_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__or3_4
Xfanout159 _04913_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout384_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ top.a1.instruction\[7\] top.a1.instruction\[8\] net745 vssd1 vssd1 vccd1
+ vccd1 _04738_ sky130_fd_sc_hd__o21a_1
X_06936_ top.DUT.register\[8\]\[22\] net593 net716 top.DUT.register\[9\]\[22\] _02052_
+ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a221o_1
XANTENNA__11303__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _01420_ net872 _04675_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__o21a_1
X_06867_ _01962_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout551_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08606_ net471 _03700_ _03708_ _02522_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout649_A _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_09586_ net916 top.pc\[27\] _04603_ _04613_ net911 vssd1 vssd1 vccd1 vccd1 _00108_
+ sky130_fd_sc_hd__o221a_1
X_06798_ top.DUT.register\[6\]\[30\] net598 net591 top.DUT.register\[20\]\[30\] _01914_
+ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ net472 net305 _03636_ _02797_ net396 vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__o32a_1
XFILLER_0_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_A _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08468_ _02833_ _03576_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ top.DUT.register\[5\]\[5\] net542 net649 top.DUT.register\[12\]\[5\] _02535_
+ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10627__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ net476 _02840_ _02839_ net396 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ net1476 net235 net511 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10361_ net2245 net244 net432 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
X_12100_ _05953_ _05955_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__or3_1
XANTENNA__07994__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ clknet_leaf_33_clk _00626_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ net1375 net254 net524 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12031_ _05885_ _05887_ _05891_ _05867_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a31o_4
XANTENNA__09735__A1 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 top.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10362__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 top.DUT.register\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07210__A2 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_4
Xfanout671 net672 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_4
Xfanout682 _01675_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_8
X_12933_ clknet_leaf_40_clk _00479_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11046__X _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09171__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12864_ clknet_leaf_12_clk _00410_ net967 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11815_ _05605_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__and2_1
X_12795_ clknet_leaf_1_clk _00341_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11746_ _05568_ _05598_ _05602_ _05603_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_32_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07277__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _05520_ _05525_ _05530_ _05533_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10537__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13416_ clknet_leaf_26_clk _00962_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net233 net1869 net376 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11270__A_N net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13347_ clknet_leaf_35_clk _00893_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10559_ net249 net1566 net504 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13278_ clknet_leaf_40_clk _00824_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12229_ net1959 net867 net832 _05687_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_102_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09346__B _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07201__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07770_ top.DUT.register\[6\]\[30\] net578 net575 top.DUT.register\[7\]\[30\] _02886_
+ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__a221o_1
X_06721_ top.DUT.register\[31\]\[3\] net669 net550 top.DUT.register\[4\]\[3\] _01837_
+ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09440_ net842 _02564_ net618 vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06652_ top.DUT.register\[20\]\[2\] net561 net644 top.DUT.register\[10\]\[2\] _01768_
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_111_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09371_ net856 _01805_ _04409_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a21o_2
X_06583_ top.DUT.register\[10\]\[0\] net644 net640 top.DUT.register\[9\]\[0\] _01697_
+ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a221o_1
XANTENNA__06992__Y _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ _03434_ _03435_ net293 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08465__B2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08253_ net477 _03280_ _03279_ net397 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10447__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout132_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ top.DUT.register\[25\]\[10\] net711 net748 top.DUT.register\[1\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08184_ net325 _02244_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06226__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06228__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07135_ top.DUT.register\[20\]\[13\] net588 net707 top.DUT.register\[7\]\[13\] _02251_
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a221o_1
XANTENNA__09965__A1 _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1041_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07066_ top.DUT.register\[27\]\[16\] net770 net754 top.DUT.register\[18\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10182__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A _01560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ top.DUT.register\[1\]\[18\] net703 net540 top.DUT.register\[5\]\[18\] _03084_
+ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a221o_1
XANTENNA__10910__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06919_ top.DUT.register\[29\]\[23\] net784 net752 top.DUT.register\[17\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a22o_1
X_09707_ _04210_ _04211_ net822 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07899_ top.DUT.register\[21\]\[24\] net571 net629 top.DUT.register\[29\]\[24\] _03015_
+ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ top.pc\[31\] _04649_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_143_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09569_ top.pc\[27\] _04590_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _05421_ _05425_ _05451_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07259__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12580_ clknet_leaf_28_clk _00126_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_176_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ _05349_ _05390_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10357__S net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
X_11462_ _05291_ _05318_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__xor2_4
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09405__B1 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire368 _01591_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
X_13201_ clknet_leaf_7_clk _00747_ net970 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10413_ net1873 net163 net515 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA__09956__A1 _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11393_ _05252_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07967__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13132_ clknet_leaf_2_clk _00678_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10344_ net1818 net177 net518 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
X_13063_ clknet_leaf_53_clk _00609_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10092__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ net185 net1402 net435 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _05846_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10820__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net492 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_4
XANTENNA__09341__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12916_ clknet_leaf_99_clk _00462_ net1004 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08695__B2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ clknet_leaf_24_clk _00393_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ clknet_leaf_2_clk _00324_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11729_ top.a1.dataIn\[9\] _05589_ _05588_ _05587_ vssd1 vssd1 vccd1 vccd1 _05590_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10267__S net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__B _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold905 top.DUT.register\[6\]\[18\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 top.DUT.register\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07958__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 top.DUT.register\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07422__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold938 top.DUT.register\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 top.DUT.register\[5\]\[0\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ _03983_ _04027_ net317 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ _03930_ _03961_ _03054_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_209_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08383__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ top.DUT.register\[22\]\[28\] net553 net656 top.DUT.register\[28\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a22o_1
XANTENNA__10730__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__A1_N _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ top.DUT.register\[19\]\[31\] net674 net669 top.DUT.register\[31\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08135__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ top.DUT.register\[28\]\[4\] net657 net637 top.DUT.register\[25\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a22o_1
X_07684_ top.DUT.register\[30\]\[12\] net695 net643 top.DUT.register\[10\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07489__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ net854 _02564_ net618 _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__o22a_4
XANTENNA__09820__A _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06635_ top.a1.instruction\[23\] _01616_ _01640_ top.a1.instruction\[31\] vssd1 vssd1
+ vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
XANTENNA__06697__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _04376_ _04379_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1089_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06566_ net747 _01652_ _01656_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__and3_1
XANTENNA__08438__B2 _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ net397 _02844_ net464 _03419_ _03416_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08989__A2 _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _04311_ _04314_ _04312_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10177__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06497_ _01512_ _01612_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ net319 net356 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07661__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09938__A1 _04622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ _02562_ _02838_ _02841_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ top.DUT.register\[10\]\[14\] net727 net719 top.DUT.register\[26\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XANTENNA__07413__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08098_ top.DUT.register\[22\]\[22\] net553 net664 top.DUT.register\[14\]\[22\] _03214_
+ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout883_A _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07058__Y _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ _02161_ _02162_ _02164_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__or4_1
X_10060_ net224 top.DUT.register\[4\]\[10\] net446 vssd1 vssd1 vccd1 vccd1 _00228_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08126__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Left_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09323__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ clknet_leaf_64_clk _01275_ net1098 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ net1724 net216 net481 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_178_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ clknet_leaf_118_clk _00247_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13681_ clknet_leaf_88_clk _01222_ net1017 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
X_10893_ net2034 net231 net408 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ clknet_leaf_36_clk _00178_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08429__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12225__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11043__Y _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10087__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ clknet_leaf_87_clk _00109_ net1016 vssd1 vssd1 vccd1 vccd1 top.pc\[28\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_81_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08065__B _03178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _05369_ _05373_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_156_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ clknet_leaf_89_clk _00041_ net1013 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06860__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ top.a1.dataIn\[17\] _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__or3_2
XANTENNA__10815__S net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11376_ top.a1.dataIn\[22\] top.a1.dataIn\[21\] top.a1.dataIn\[20\] vssd1 vssd1 vccd1
+ vccd1 _05237_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_189_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10327_ net2205 net251 net519 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ clknet_leaf_5_clk _00661_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_13046_ clknet_leaf_102_clk _00592_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09905__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ net267 net2037 net437 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__mux2_1
XANTENNA__10550__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ net257 top.DUT.register\[8\]\[2\] net439 vssd1 vssd1 vccd1 vccd1 _00348_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13879_ net1139 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_201_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06420_ net810 _01535_ _01536_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and3_1
XANTENNA__07431__Y _02548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06351_ _01335_ _01468_ _01478_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09070_ _04116_ _04119_ _04120_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or4_1
XFILLER_0_142_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06282_ net2239 net898 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[8\] sky130_fd_sc_hd__and2_1
XFILLER_0_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07643__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__B2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08021_ top.DUT.register\[26\]\[19\] net679 net659 top.DUT.register\[18\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06851__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10725__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13652__CLK clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 top.DUT.register\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09087__A _03927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09396__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold713 top.DUT.register\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold724 top.DUT.register\[8\]\[0\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold735 top.DUT.register\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold746 top.DUT.register\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 top.DUT.register\[12\]\[29\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__B1 _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold768 top.DUT.register\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold779 top.DUT.register\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _04669_ net361 net329 top.a1.dataIn\[31\] net364 vssd1 vssd1 vccd1 vccd1
+ _04955_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08923_ _03963_ _04011_ _03005_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10460__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net275 _03378_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1004_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ top.DUT.register\[26\]\[29\] net679 net675 top.DUT.register\[13\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ net1304 net859 net837 _03880_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a22o_1
XANTENNA__08108__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout464_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07736_ _02694_ _02745_ _02799_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__or4_1
XFILLER_0_211_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09856__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ top.DUT.register\[6\]\[10\] net576 net683 top.DUT.register\[2\]\[10\] _02783_
+ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout631_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__Y _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06618_ _01599_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__or2_4
X_09406_ net841 _01803_ net619 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21oi_1
X_07598_ net829 _02714_ net468 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07882__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _02264_ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__or2_1
X_06549_ net747 _01649_ _01653_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06425__A_N top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _02346_ _02668_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__nor2_1
XANTENNA__07634__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ net299 _02109_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__and2_1
XANTENNA__06842__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09199_ _04232_ _04235_ _04248_ _01632_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o31a_1
XANTENNA__10635__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11230_ _05115_ net1302 net402 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07398__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ net922 net1346 net874 _05080_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a31o_1
X_10112_ net150 net2081 net387 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__mux2_1
X_11092_ net1198 net878 net846 top.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 _01171_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ net148 net2098 net529 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
XANTENNA__10370__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__A1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 _01178_ vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__B2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 top.lcd.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _01170_ vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 _01180_ vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold84 net97 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 top.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_69_clk _01327_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11994_ _05821_ _05833_ _05810_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09460__A _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_62_clk _01263_ net1108 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ net2090 net152 net487 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13664_ clknet_leaf_90_clk _01205_ net1003 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
X_10876_ net2196 net165 net491 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
XANTENNA__07873__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12615_ clknet_leaf_44_clk _00161_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13595_ clknet_leaf_55_clk _01136_ net1093 vssd1 vssd1 vccd1 vccd1 top.ramload\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12546_ clknet_leaf_98_clk _00092_ net1005 vssd1 vssd1 vccd1 vccd1 top.pc\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06833__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10545__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__B _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ clknet_leaf_87_clk _00024_ net1017 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_4 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ _05261_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11359_ top.a1.dataIn\[23\] _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08050__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10280__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13029_ clknet_leaf_47_clk _00575_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08889__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1073 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_2
XANTENNA__07010__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1084 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1095 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
XANTENNA__13117__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08570_ net311 _03674_ _03673_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07521_ net825 _02637_ _02617_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07452_ top.DUT.register\[11\]\[6\] net702 net555 top.DUT.register\[22\]\[6\] _02568_
+ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06403_ top.a1.instruction\[18\] _01519_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11124__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ top.DUT.register\[9\]\[4\] net718 net753 top.DUT.register\[17\]\[4\] _02499_
+ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09122_ top.a1.instruction\[12\] _01604_ _01498_ vssd1 vssd1 vccd1 vccd1 _04175_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06334_ _01462_ _01463_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a22o_1
XANTENNA__07616__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _03642_ _03651_ _03693_ _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__and4_1
XFILLER_0_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10455__S net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06265_ net1241 net892 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[23\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08004_ top.DUT.register\[2\]\[21\] net684 net644 top.DUT.register\[10\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__a22o_1
Xhold510 top.DUT.register\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06196_ top.pc\[31\] vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
Xhold521 top.DUT.register\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 top.DUT.register\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 top.DUT.register\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 top.pad.keyCode\[3\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 top.DUT.register\[16\]\[1\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1121_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 top.lcd.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 top.DUT.register\[22\]\[18\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 top.DUT.register\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _04938_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout581_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_A _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10190__S net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _03978_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__and2b_1
X_09886_ _03897_ net455 net534 _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout1007_X net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1210 top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08837_ _03180_ _03914_ _03032_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _03082_ _03840_ _03081_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07719_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ _02519_ _03786_ _03798_ net466 _03796_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ net222 net1584 net415 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XANTENNA__07855__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ net234 net1636 net420 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ clknet_leaf_60_clk _00008_ net1102 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07068__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13380_ clknet_leaf_29_clk _00926_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ net252 net1745 net424 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07607__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12422__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ top.lcd.cnt_500hz\[12\] _06123_ net743 vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_153_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06815__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__S net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ _06080_ _06083_ net1119 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11213_ net1257 net404 net369 _05109_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_186_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12193_ _06044_ _06047_ _06048_ _06045_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a22oi_2
XANTENNA__08032__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_208_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11144_ net46 net882 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__and2_1
XANTENNA__07240__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A2 _04198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ net22 net863 net835 net1382 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__o22a_1
X_10026_ net216 net1756 net529 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XANTENNA_input28_X net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_201_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08099__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11977_ _05802_ _05834_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13716_ clknet_leaf_65_clk _01246_ net1112 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ net1681 net221 net486 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__mux2_1
XANTENNA__07846__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ clknet_leaf_93_clk net1230 net995 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
X_10859_ net1553 net235 net491 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08694__A1_N net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13578_ clknet_leaf_55_clk _01119_ net1097 vssd1 vssd1 vccd1 vccd1 top.a1.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_167_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06806__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ clknet_leaf_44_clk _00075_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10275__S net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08023__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net312 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_0_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09740_ net265 net1738 net393 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__mux2_1
X_06952_ net325 _02068_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nand2_1
.ends

