VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO team_12_Wrapper
  CLASS BLOCK ;
  FOREIGN team_12_Wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 899.000 ;
  PIN ACK_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END ACK_I
  PIN ADR_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END ADR_O[0]
  PIN ADR_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END ADR_O[10]
  PIN ADR_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END ADR_O[11]
  PIN ADR_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END ADR_O[12]
  PIN ADR_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END ADR_O[13]
  PIN ADR_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END ADR_O[14]
  PIN ADR_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END ADR_O[15]
  PIN ADR_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END ADR_O[16]
  PIN ADR_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END ADR_O[17]
  PIN ADR_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END ADR_O[18]
  PIN ADR_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END ADR_O[19]
  PIN ADR_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END ADR_O[1]
  PIN ADR_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END ADR_O[20]
  PIN ADR_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END ADR_O[21]
  PIN ADR_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 574.640 800.000 575.240 ;
    END
  END ADR_O[22]
  PIN ADR_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 391.040 800.000 391.640 ;
    END
  END ADR_O[23]
  PIN ADR_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 448.840 800.000 449.440 ;
    END
  END ADR_O[24]
  PIN ADR_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.040 800.000 425.640 ;
    END
  END ADR_O[25]
  PIN ADR_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END ADR_O[26]
  PIN ADR_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END ADR_O[27]
  PIN ADR_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END ADR_O[28]
  PIN ADR_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END ADR_O[29]
  PIN ADR_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END ADR_O[2]
  PIN ADR_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END ADR_O[30]
  PIN ADR_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 591.640 800.000 592.240 ;
    END
  END ADR_O[31]
  PIN ADR_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END ADR_O[3]
  PIN ADR_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END ADR_O[4]
  PIN ADR_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 482.840 800.000 483.440 ;
    END
  END ADR_O[5]
  PIN ADR_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END ADR_O[6]
  PIN ADR_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END ADR_O[7]
  PIN ADR_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END ADR_O[8]
  PIN ADR_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END ADR_O[9]
  PIN CYC_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 527.040 800.000 527.640 ;
    END
  END CYC_O
  PIN DAT_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END DAT_I[0]
  PIN DAT_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END DAT_I[10]
  PIN DAT_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END DAT_I[11]
  PIN DAT_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END DAT_I[12]
  PIN DAT_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END DAT_I[13]
  PIN DAT_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END DAT_I[14]
  PIN DAT_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END DAT_I[15]
  PIN DAT_I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END DAT_I[16]
  PIN DAT_I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END DAT_I[17]
  PIN DAT_I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END DAT_I[18]
  PIN DAT_I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END DAT_I[19]
  PIN DAT_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END DAT_I[1]
  PIN DAT_I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END DAT_I[20]
  PIN DAT_I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END DAT_I[21]
  PIN DAT_I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END DAT_I[22]
  PIN DAT_I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END DAT_I[23]
  PIN DAT_I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END DAT_I[24]
  PIN DAT_I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END DAT_I[25]
  PIN DAT_I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END DAT_I[26]
  PIN DAT_I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END DAT_I[27]
  PIN DAT_I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END DAT_I[28]
  PIN DAT_I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END DAT_I[29]
  PIN DAT_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END DAT_I[2]
  PIN DAT_I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END DAT_I[30]
  PIN DAT_I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END DAT_I[31]
  PIN DAT_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END DAT_I[3]
  PIN DAT_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END DAT_I[4]
  PIN DAT_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END DAT_I[5]
  PIN DAT_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END DAT_I[6]
  PIN DAT_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END DAT_I[7]
  PIN DAT_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END DAT_I[8]
  PIN DAT_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END DAT_I[9]
  PIN DAT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 261.840 800.000 262.440 ;
    END
  END DAT_O[0]
  PIN DAT_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END DAT_O[10]
  PIN DAT_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END DAT_O[11]
  PIN DAT_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 367.240 800.000 367.840 ;
    END
  END DAT_O[12]
  PIN DAT_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END DAT_O[13]
  PIN DAT_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END DAT_O[14]
  PIN DAT_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END DAT_O[15]
  PIN DAT_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END DAT_O[16]
  PIN DAT_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 397.840 800.000 398.440 ;
    END
  END DAT_O[17]
  PIN DAT_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END DAT_O[18]
  PIN DAT_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END DAT_O[19]
  PIN DAT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END DAT_O[1]
  PIN DAT_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END DAT_O[20]
  PIN DAT_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END DAT_O[21]
  PIN DAT_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END DAT_O[22]
  PIN DAT_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END DAT_O[23]
  PIN DAT_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END DAT_O[24]
  PIN DAT_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END DAT_O[25]
  PIN DAT_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END DAT_O[26]
  PIN DAT_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END DAT_O[27]
  PIN DAT_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END DAT_O[28]
  PIN DAT_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END DAT_O[29]
  PIN DAT_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END DAT_O[2]
  PIN DAT_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END DAT_O[30]
  PIN DAT_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END DAT_O[31]
  PIN DAT_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 224.440 800.000 225.040 ;
    END
  END DAT_O[3]
  PIN DAT_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 374.040 800.000 374.640 ;
    END
  END DAT_O[4]
  PIN DAT_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 547.440 800.000 548.040 ;
    END
  END DAT_O[5]
  PIN DAT_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END DAT_O[6]
  PIN DAT_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 173.440 800.000 174.040 ;
    END
  END DAT_O[7]
  PIN DAT_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 91.840 800.000 92.440 ;
    END
  END DAT_O[8]
  PIN DAT_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 23.840 800.000 24.440 ;
    END
  END DAT_O[9]
  PIN SEL_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 469.240 800.000 469.840 ;
    END
  END SEL_O[0]
  PIN SEL_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 190.440 800.000 191.040 ;
    END
  END SEL_O[1]
  PIN SEL_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 214.240 800.000 214.840 ;
    END
  END SEL_O[2]
  PIN SEL_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 588.240 800.000 588.840 ;
    END
  END SEL_O[3]
  PIN STB_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 578.040 800.000 578.640 ;
    END
  END STB_O
  PIN WE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 221.040 800.000 221.640 ;
    END
  END WE_O
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 154.650 895.000 154.930 899.000 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END gpio_in[33]
  PIN gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END gpio_in[34]
  PIN gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END gpio_in[35]
  PIN gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END gpio_in[36]
  PIN gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END gpio_in[37]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 796.000 741.240 800.000 741.840 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END gpio_in[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 890.840 800.000 891.440 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 499.840 800.000 500.440 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 608.640 800.000 609.240 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 88.440 800.000 89.040 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 581.440 800.000 582.040 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 149.640 800.000 150.240 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 159.840 800.000 160.440 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 544.040 800.000 544.640 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 146.240 800.000 146.840 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 401.240 800.000 401.840 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 136.040 800.000 136.640 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 880.640 800.000 881.240 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 295.840 800.000 296.440 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 513.440 800.000 514.040 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 139.440 800.000 140.040 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 6.840 800.000 7.440 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 156.440 800.000 157.040 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 438.640 800.000 439.240 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 472.640 800.000 473.240 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 363.840 800.000 364.440 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 489.640 800.000 490.240 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 404.640 800.000 405.240 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 877.240 800.000 877.840 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 462.440 800.000 463.040 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 193.840 800.000 194.440 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 47.640 800.000 48.240 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 567.840 800.000 568.440 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.240 800.000 350.840 ;
    END
  END gpio_oeb[34]
  PIN gpio_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 459.040 800.000 459.640 ;
    END
  END gpio_oeb[35]
  PIN gpio_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 377.440 800.000 378.040 ;
    END
  END gpio_oeb[36]
  PIN gpio_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 625.640 800.000 626.240 ;
    END
  END gpio_oeb[37]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 873.840 800.000 874.440 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 887.440 800.000 888.040 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 884.040 800.000 884.640 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 870.440 800.000 871.040 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.240 800.000 299.840 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 85.040 800.000 85.640 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 340.040 800.000 340.640 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 122.440 800.000 123.040 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 724.240 800.000 724.840 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 693.640 800.000 694.240 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 683.440 800.000 684.040 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 697.040 800.000 697.640 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 717.440 800.000 718.040 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 727.640 800.000 728.240 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 690.240 800.000 690.840 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 731.040 800.000 731.640 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 700.440 800.000 701.040 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 680.040 800.000 680.640 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 115.640 800.000 116.240 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 707.240 800.000 707.840 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 720.840 800.000 721.440 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 734.440 800.000 735.040 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 258.440 800.000 259.040 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 323.040 800.000 323.640 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 455.640 800.000 456.240 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 78.240 800.000 78.840 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 170.040 800.000 170.640 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 17.040 800.000 17.640 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 428.440 800.000 429.040 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 309.440 800.000 310.040 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.240 800.000 316.840 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 153.040 800.000 153.640 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 336.640 800.000 337.240 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 0.040 800.000 0.640 ;
    END
  END gpio_out[33]
  PIN gpio_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 30.640 800.000 31.240 ;
    END
  END gpio_out[34]
  PIN gpio_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 57.840 800.000 58.440 ;
    END
  END gpio_out[35]
  PIN gpio_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 95.240 800.000 95.840 ;
    END
  END gpio_out[36]
  PIN gpio_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 329.840 800.000 330.440 ;
    END
  END gpio_out[37]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 418.240 800.000 418.840 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 71.440 800.000 72.040 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 659.640 800.000 660.240 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 282.240 800.000 282.840 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 710.640 800.000 711.240 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 737.840 800.000 738.440 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 714.040 800.000 714.640 ;
    END
  END gpio_out[9]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 408.040 800.000 408.640 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 200.640 800.000 201.240 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 486.240 800.000 486.840 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 40.840 800.000 41.440 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 265.240 800.000 265.840 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 605.240 800.000 605.840 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 119.040 800.000 119.640 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 241.440 800.000 242.040 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 652.840 800.000 653.440 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.240 800.000 384.840 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 61.240 800.000 61.840 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 217.640 800.000 218.240 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 68.040 800.000 68.640 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 629.040 800.000 629.640 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 231.240 800.000 231.840 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 479.440 800.000 480.040 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 272.040 800.000 272.640 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 255.040 800.000 255.640 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 125.840 800.000 126.440 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 476.040 800.000 476.640 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 571.240 800.000 571.840 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 506.640 800.000 507.240 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 10.240 800.000 10.840 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 414.840 800.000 415.440 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 431.840 800.000 432.440 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 238.040 800.000 238.640 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 98.640 800.000 99.240 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 520.240 800.000 520.840 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 142.840 800.000 143.440 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 646.040 800.000 646.640 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 204.040 800.000 204.640 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 278.840 800.000 279.440 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 289.040 800.000 289.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 380.840 800.000 381.440 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 584.840 800.000 585.440 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 465.840 800.000 466.440 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 649.440 800.000 650.040 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 333.240 800.000 333.840 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 180.240 800.000 180.840 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 676.640 800.000 677.240 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 37.440 800.000 38.040 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 435.240 800.000 435.840 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 112.240 800.000 112.840 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 248.240 800.000 248.840 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 530.440 800.000 531.040 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 34.040 800.000 34.640 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 622.240 800.000 622.840 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 442.040 800.000 442.640 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 595.040 800.000 595.640 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 105.440 800.000 106.040 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 360.440 800.000 361.040 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 635.840 800.000 636.440 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 523.640 800.000 524.240 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 108.840 800.000 109.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 550.840 800.000 551.440 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.040 800.000 51.640 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 618.840 800.000 619.440 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 540.640 800.000 541.240 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 663.040 800.000 663.640 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 302.640 800.000 303.240 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 183.640 800.000 184.240 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 27.240 800.000 27.840 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 357.040 800.000 357.640 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 666.440 800.000 667.040 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 642.640 800.000 643.240 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 346.840 800.000 347.440 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 3.440 800.000 4.040 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 353.640 800.000 354.240 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 20.440 800.000 21.040 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 268.640 800.000 269.240 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 533.840 800.000 534.440 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 615.440 800.000 616.040 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 510.040 800.000 510.640 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 285.640 800.000 286.240 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 639.240 800.000 639.840 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 244.840 800.000 245.440 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 306.040 800.000 306.640 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 251.640 800.000 252.240 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 54.440 800.000 55.040 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 669.840 800.000 670.440 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 601.840 800.000 602.440 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 163.240 800.000 163.840 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 312.840 800.000 313.440 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 227.840 800.000 228.440 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 421.640 800.000 422.240 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 187.040 800.000 187.640 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 673.240 800.000 673.840 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 132.640 800.000 133.240 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 370.640 800.000 371.240 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.040 800.000 493.640 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 13.640 800.000 14.240 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 197.240 800.000 197.840 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 656.240 800.000 656.840 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 561.040 800.000 561.640 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 503.240 800.000 503.840 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 554.240 800.000 554.840 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 234.640 800.000 235.240 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 81.640 800.000 82.240 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 44.240 800.000 44.840 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 557.640 800.000 558.240 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 387.640 800.000 388.240 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 632.440 800.000 633.040 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 102.040 800.000 102.640 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 319.640 800.000 320.240 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 496.440 800.000 497.040 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 516.840 800.000 517.440 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 129.240 800.000 129.840 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 166.640 800.000 167.240 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 292.440 800.000 293.040 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 64.640 800.000 65.240 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 275.440 800.000 276.040 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 612.040 800.000 612.640 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 598.440 800.000 599.040 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 394.440 800.000 395.040 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 564.440 800.000 565.040 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 343.440 800.000 344.040 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 74.840 800.000 75.440 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 326.440 800.000 327.040 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 207.440 800.000 208.040 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 452.240 800.000 452.840 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 537.240 800.000 537.840 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 411.440 800.000 412.040 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 445.440 800.000 446.040 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 703.840 800.000 704.440 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 686.840 800.000 687.440 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 894.240 800.000 894.840 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 744.640 800.000 745.240 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 897.640 800.000 898.240 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 748.040 800.000 748.640 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 751.440 800.000 752.040 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 754.840 800.000 755.440 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 758.240 800.000 758.840 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 761.640 800.000 762.240 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 765.040 800.000 765.640 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 768.440 800.000 769.040 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 771.840 800.000 772.440 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 775.240 800.000 775.840 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 778.640 800.000 779.240 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 782.040 800.000 782.640 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 785.440 800.000 786.040 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 788.840 800.000 789.440 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 792.240 800.000 792.840 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 795.640 800.000 796.240 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 799.040 800.000 799.640 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 802.440 800.000 803.040 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 805.840 800.000 806.440 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 809.240 800.000 809.840 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 812.640 800.000 813.240 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 816.040 800.000 816.640 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 819.440 800.000 820.040 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 822.840 800.000 823.440 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 826.240 800.000 826.840 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 829.640 800.000 830.240 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 833.040 800.000 833.640 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 836.440 800.000 837.040 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 839.840 800.000 840.440 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 843.240 800.000 843.840 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 846.640 800.000 847.240 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 850.040 800.000 850.640 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 853.440 800.000 854.040 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 856.840 800.000 857.440 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 860.240 800.000 860.840 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 863.640 800.000 864.240 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 867.040 800.000 867.640 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 895.000 798.930 899.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 895.000 795.710 899.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 895.000 792.490 899.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 895.000 789.270 899.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 895.000 786.050 899.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 895.000 782.830 899.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 895.000 779.610 899.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 895.000 776.390 899.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 895.000 773.170 899.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 895.000 769.950 899.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 895.000 766.730 899.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 895.000 763.510 899.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 895.000 760.290 899.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 895.000 757.070 899.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 895.000 753.850 899.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 895.000 750.630 899.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 895.000 747.410 899.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 895.000 744.190 899.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 895.000 740.970 899.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 895.000 737.750 899.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 895.000 734.530 899.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 895.000 731.310 899.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 895.000 728.090 899.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 895.000 724.870 899.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 895.000 721.650 899.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 895.000 718.430 899.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 895.000 715.210 899.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 895.000 711.990 899.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 895.000 708.770 899.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 895.000 705.550 899.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 895.000 702.330 899.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 895.000 699.110 899.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 895.000 695.890 899.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 895.000 692.670 899.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 895.000 689.450 899.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 895.000 686.230 899.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 895.000 683.010 899.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 895.000 679.790 899.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 895.000 676.570 899.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 895.000 673.350 899.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 895.000 670.130 899.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 895.000 666.910 899.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 895.000 663.690 899.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 895.000 660.470 899.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 895.000 657.250 899.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 895.000 654.030 899.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 895.000 650.810 899.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 895.000 647.590 899.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 895.000 644.370 899.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 895.000 641.150 899.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 895.000 637.930 899.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 895.000 634.710 899.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 895.000 631.490 899.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 895.000 628.270 899.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 895.000 625.050 899.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 895.000 621.830 899.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 895.000 618.610 899.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 895.000 615.390 899.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 895.000 612.170 899.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 895.000 608.950 899.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 895.000 605.730 899.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 895.000 602.510 899.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 895.000 599.290 899.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 895.000 596.070 899.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 895.000 592.850 899.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 895.000 589.630 899.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 895.000 586.410 899.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 895.000 583.190 899.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 895.000 579.970 899.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 895.000 576.750 899.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 895.000 573.530 899.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 895.000 570.310 899.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 895.000 567.090 899.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 895.000 563.870 899.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 895.000 560.650 899.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 895.000 557.430 899.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 895.000 554.210 899.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 895.000 550.990 899.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 895.000 547.770 899.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 895.000 544.550 899.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 895.000 541.330 899.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 895.000 538.110 899.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 895.000 534.890 899.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 895.000 531.670 899.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 895.000 528.450 899.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 895.000 525.230 899.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 895.000 522.010 899.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 895.000 518.790 899.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 895.000 515.570 899.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 886.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 895.000 16.470 899.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 61.270 895.000 61.550 899.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.970 895.000 13.250 899.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 895.000 45.450 899.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.050 895.000 58.330 899.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 96.690 895.000 96.970 899.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 895.000 77.650 899.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 895.000 32.570 899.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 25.850 895.000 26.130 899.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 125.670 895.000 125.950 899.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 895.000 29.350 899.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 895.000 109.850 899.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.950 895.000 42.230 899.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 3.310 895.000 3.590 899.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.550 895.000 138.830 899.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 0.090 895.000 0.370 899.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.750 895.000 10.030 899.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 895.000 39.010 899.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 895.000 116.290 899.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 895.000 145.270 899.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.770 895.000 142.050 899.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.530 895.000 6.810 899.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 895.000 135.610 899.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 895.000 90.530 899.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 895.000 19.690 899.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 895.000 51.890 899.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.930 895.000 71.210 899.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.910 895.000 100.190 899.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.150 895.000 74.430 899.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.510 895.000 35.790 899.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.830 895.000 55.110 899.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 119.230 895.000 119.510 899.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.710 895.000 67.990 899.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.790 895.000 113.070 899.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.130 895.000 103.410 899.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 895.000 512.350 899.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 895.000 509.130 899.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 895.000 505.910 899.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 895.000 502.690 899.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 895.000 499.470 899.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 895.000 496.250 899.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 895.000 493.030 899.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 895.000 489.810 899.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 895.000 486.590 899.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 895.000 483.370 899.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 895.000 480.150 899.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 895.000 476.930 899.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 895.000 473.710 899.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 895.000 470.490 899.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 895.000 467.270 899.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 895.000 464.050 899.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 895.000 460.830 899.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 895.000 457.610 899.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 895.000 454.390 899.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 895.000 451.170 899.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 895.000 447.950 899.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 895.000 444.730 899.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 895.000 441.510 899.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 895.000 438.290 899.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 895.000 435.070 899.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 895.000 431.850 899.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 895.000 428.630 899.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 895.000 425.410 899.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 895.000 422.190 899.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 895.000 418.970 899.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 895.000 415.750 899.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 895.000 93.750 899.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 895.000 106.630 899.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 128.890 895.000 129.170 899.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 895.000 22.910 899.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 895.000 84.090 899.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 895.000 80.870 899.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 895.000 151.710 899.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 895.000 132.390 899.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 895.000 48.670 899.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 895.000 122.730 899.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 895.000 87.310 899.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 895.000 64.770 899.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.210 895.000 148.490 899.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 895.000 412.530 899.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 895.000 409.310 899.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 895.000 406.090 899.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 895.000 402.870 899.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 886.805 ;
      LAYER met1 ;
        RECT 0.070 10.640 798.950 889.740 ;
      LAYER met2 ;
        RECT 0.650 894.720 3.030 895.290 ;
        RECT 3.870 894.720 6.250 895.290 ;
        RECT 7.090 894.720 9.470 895.290 ;
        RECT 10.310 894.720 12.690 895.290 ;
        RECT 13.530 894.720 15.910 895.290 ;
        RECT 16.750 894.720 19.130 895.290 ;
        RECT 19.970 894.720 22.350 895.290 ;
        RECT 23.190 894.720 25.570 895.290 ;
        RECT 26.410 894.720 28.790 895.290 ;
        RECT 29.630 894.720 32.010 895.290 ;
        RECT 32.850 894.720 35.230 895.290 ;
        RECT 36.070 894.720 38.450 895.290 ;
        RECT 39.290 894.720 41.670 895.290 ;
        RECT 42.510 894.720 44.890 895.290 ;
        RECT 45.730 894.720 48.110 895.290 ;
        RECT 48.950 894.720 51.330 895.290 ;
        RECT 52.170 894.720 54.550 895.290 ;
        RECT 55.390 894.720 57.770 895.290 ;
        RECT 58.610 894.720 60.990 895.290 ;
        RECT 61.830 894.720 64.210 895.290 ;
        RECT 65.050 894.720 67.430 895.290 ;
        RECT 68.270 894.720 70.650 895.290 ;
        RECT 71.490 894.720 73.870 895.290 ;
        RECT 74.710 894.720 77.090 895.290 ;
        RECT 77.930 894.720 80.310 895.290 ;
        RECT 81.150 894.720 83.530 895.290 ;
        RECT 84.370 894.720 86.750 895.290 ;
        RECT 87.590 894.720 89.970 895.290 ;
        RECT 90.810 894.720 93.190 895.290 ;
        RECT 94.030 894.720 96.410 895.290 ;
        RECT 97.250 894.720 99.630 895.290 ;
        RECT 100.470 894.720 102.850 895.290 ;
        RECT 103.690 894.720 106.070 895.290 ;
        RECT 106.910 894.720 109.290 895.290 ;
        RECT 110.130 894.720 112.510 895.290 ;
        RECT 113.350 894.720 115.730 895.290 ;
        RECT 116.570 894.720 118.950 895.290 ;
        RECT 119.790 894.720 122.170 895.290 ;
        RECT 123.010 894.720 125.390 895.290 ;
        RECT 126.230 894.720 128.610 895.290 ;
        RECT 129.450 894.720 131.830 895.290 ;
        RECT 132.670 894.720 135.050 895.290 ;
        RECT 135.890 894.720 138.270 895.290 ;
        RECT 139.110 894.720 141.490 895.290 ;
        RECT 142.330 894.720 144.710 895.290 ;
        RECT 145.550 894.720 147.930 895.290 ;
        RECT 148.770 894.720 151.150 895.290 ;
        RECT 151.990 894.720 154.370 895.290 ;
        RECT 155.210 894.720 402.310 895.290 ;
        RECT 403.150 894.720 405.530 895.290 ;
        RECT 406.370 894.720 408.750 895.290 ;
        RECT 409.590 894.720 411.970 895.290 ;
        RECT 412.810 894.720 415.190 895.290 ;
        RECT 416.030 894.720 418.410 895.290 ;
        RECT 419.250 894.720 421.630 895.290 ;
        RECT 422.470 894.720 424.850 895.290 ;
        RECT 425.690 894.720 428.070 895.290 ;
        RECT 428.910 894.720 431.290 895.290 ;
        RECT 432.130 894.720 434.510 895.290 ;
        RECT 435.350 894.720 437.730 895.290 ;
        RECT 438.570 894.720 440.950 895.290 ;
        RECT 441.790 894.720 444.170 895.290 ;
        RECT 445.010 894.720 447.390 895.290 ;
        RECT 448.230 894.720 450.610 895.290 ;
        RECT 451.450 894.720 453.830 895.290 ;
        RECT 454.670 894.720 457.050 895.290 ;
        RECT 457.890 894.720 460.270 895.290 ;
        RECT 461.110 894.720 463.490 895.290 ;
        RECT 464.330 894.720 466.710 895.290 ;
        RECT 467.550 894.720 469.930 895.290 ;
        RECT 470.770 894.720 473.150 895.290 ;
        RECT 473.990 894.720 476.370 895.290 ;
        RECT 477.210 894.720 479.590 895.290 ;
        RECT 480.430 894.720 482.810 895.290 ;
        RECT 483.650 894.720 486.030 895.290 ;
        RECT 486.870 894.720 489.250 895.290 ;
        RECT 490.090 894.720 492.470 895.290 ;
        RECT 493.310 894.720 495.690 895.290 ;
        RECT 496.530 894.720 498.910 895.290 ;
        RECT 499.750 894.720 502.130 895.290 ;
        RECT 502.970 894.720 505.350 895.290 ;
        RECT 506.190 894.720 508.570 895.290 ;
        RECT 509.410 894.720 511.790 895.290 ;
        RECT 512.630 894.720 515.010 895.290 ;
        RECT 515.850 894.720 518.230 895.290 ;
        RECT 519.070 894.720 521.450 895.290 ;
        RECT 522.290 894.720 524.670 895.290 ;
        RECT 525.510 894.720 527.890 895.290 ;
        RECT 528.730 894.720 531.110 895.290 ;
        RECT 531.950 894.720 534.330 895.290 ;
        RECT 535.170 894.720 537.550 895.290 ;
        RECT 538.390 894.720 540.770 895.290 ;
        RECT 541.610 894.720 543.990 895.290 ;
        RECT 544.830 894.720 547.210 895.290 ;
        RECT 548.050 894.720 550.430 895.290 ;
        RECT 551.270 894.720 553.650 895.290 ;
        RECT 554.490 894.720 556.870 895.290 ;
        RECT 557.710 894.720 560.090 895.290 ;
        RECT 560.930 894.720 563.310 895.290 ;
        RECT 564.150 894.720 566.530 895.290 ;
        RECT 567.370 894.720 569.750 895.290 ;
        RECT 570.590 894.720 572.970 895.290 ;
        RECT 573.810 894.720 576.190 895.290 ;
        RECT 577.030 894.720 579.410 895.290 ;
        RECT 580.250 894.720 582.630 895.290 ;
        RECT 583.470 894.720 585.850 895.290 ;
        RECT 586.690 894.720 589.070 895.290 ;
        RECT 589.910 894.720 592.290 895.290 ;
        RECT 593.130 894.720 595.510 895.290 ;
        RECT 596.350 894.720 598.730 895.290 ;
        RECT 599.570 894.720 601.950 895.290 ;
        RECT 602.790 894.720 605.170 895.290 ;
        RECT 606.010 894.720 608.390 895.290 ;
        RECT 609.230 894.720 611.610 895.290 ;
        RECT 612.450 894.720 614.830 895.290 ;
        RECT 615.670 894.720 618.050 895.290 ;
        RECT 618.890 894.720 621.270 895.290 ;
        RECT 622.110 894.720 624.490 895.290 ;
        RECT 625.330 894.720 627.710 895.290 ;
        RECT 628.550 894.720 630.930 895.290 ;
        RECT 631.770 894.720 634.150 895.290 ;
        RECT 634.990 894.720 637.370 895.290 ;
        RECT 638.210 894.720 640.590 895.290 ;
        RECT 641.430 894.720 643.810 895.290 ;
        RECT 644.650 894.720 647.030 895.290 ;
        RECT 647.870 894.720 650.250 895.290 ;
        RECT 651.090 894.720 653.470 895.290 ;
        RECT 654.310 894.720 656.690 895.290 ;
        RECT 657.530 894.720 659.910 895.290 ;
        RECT 660.750 894.720 663.130 895.290 ;
        RECT 663.970 894.720 666.350 895.290 ;
        RECT 667.190 894.720 669.570 895.290 ;
        RECT 670.410 894.720 672.790 895.290 ;
        RECT 673.630 894.720 676.010 895.290 ;
        RECT 676.850 894.720 679.230 895.290 ;
        RECT 680.070 894.720 682.450 895.290 ;
        RECT 683.290 894.720 685.670 895.290 ;
        RECT 686.510 894.720 688.890 895.290 ;
        RECT 689.730 894.720 692.110 895.290 ;
        RECT 692.950 894.720 695.330 895.290 ;
        RECT 696.170 894.720 698.550 895.290 ;
        RECT 699.390 894.720 701.770 895.290 ;
        RECT 702.610 894.720 704.990 895.290 ;
        RECT 705.830 894.720 708.210 895.290 ;
        RECT 709.050 894.720 711.430 895.290 ;
        RECT 712.270 894.720 714.650 895.290 ;
        RECT 715.490 894.720 717.870 895.290 ;
        RECT 718.710 894.720 721.090 895.290 ;
        RECT 721.930 894.720 724.310 895.290 ;
        RECT 725.150 894.720 727.530 895.290 ;
        RECT 728.370 894.720 730.750 895.290 ;
        RECT 731.590 894.720 733.970 895.290 ;
        RECT 734.810 894.720 737.190 895.290 ;
        RECT 738.030 894.720 740.410 895.290 ;
        RECT 741.250 894.720 743.630 895.290 ;
        RECT 744.470 894.720 746.850 895.290 ;
        RECT 747.690 894.720 750.070 895.290 ;
        RECT 750.910 894.720 753.290 895.290 ;
        RECT 754.130 894.720 756.510 895.290 ;
        RECT 757.350 894.720 759.730 895.290 ;
        RECT 760.570 894.720 762.950 895.290 ;
        RECT 763.790 894.720 766.170 895.290 ;
        RECT 767.010 894.720 769.390 895.290 ;
        RECT 770.230 894.720 772.610 895.290 ;
        RECT 773.450 894.720 775.830 895.290 ;
        RECT 776.670 894.720 779.050 895.290 ;
        RECT 779.890 894.720 782.270 895.290 ;
        RECT 783.110 894.720 785.490 895.290 ;
        RECT 786.330 894.720 788.710 895.290 ;
        RECT 789.550 894.720 791.930 895.290 ;
        RECT 792.770 894.720 795.150 895.290 ;
        RECT 795.990 894.720 798.370 895.290 ;
        RECT 0.100 4.280 798.920 894.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.150 4.280 ;
        RECT 151.990 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 254.190 4.280 ;
        RECT 255.030 0.155 257.410 4.280 ;
        RECT 258.250 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 305.710 4.280 ;
        RECT 306.550 0.155 308.930 4.280 ;
        RECT 309.770 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 334.690 4.280 ;
        RECT 335.530 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 357.230 4.280 ;
        RECT 358.070 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 376.550 4.280 ;
        RECT 377.390 0.155 379.770 4.280 ;
        RECT 380.610 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 399.090 4.280 ;
        RECT 399.930 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 408.750 4.280 ;
        RECT 409.590 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 418.410 4.280 ;
        RECT 419.250 0.155 421.630 4.280 ;
        RECT 422.470 0.155 424.850 4.280 ;
        RECT 425.690 0.155 428.070 4.280 ;
        RECT 428.910 0.155 431.290 4.280 ;
        RECT 432.130 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 444.170 4.280 ;
        RECT 445.010 0.155 447.390 4.280 ;
        RECT 448.230 0.155 450.610 4.280 ;
        RECT 451.450 0.155 453.830 4.280 ;
        RECT 454.670 0.155 457.050 4.280 ;
        RECT 457.890 0.155 460.270 4.280 ;
        RECT 461.110 0.155 463.490 4.280 ;
        RECT 464.330 0.155 466.710 4.280 ;
        RECT 467.550 0.155 469.930 4.280 ;
        RECT 470.770 0.155 473.150 4.280 ;
        RECT 473.990 0.155 476.370 4.280 ;
        RECT 477.210 0.155 479.590 4.280 ;
        RECT 480.430 0.155 482.810 4.280 ;
        RECT 483.650 0.155 486.030 4.280 ;
        RECT 486.870 0.155 489.250 4.280 ;
        RECT 490.090 0.155 492.470 4.280 ;
        RECT 493.310 0.155 495.690 4.280 ;
        RECT 496.530 0.155 498.910 4.280 ;
        RECT 499.750 0.155 502.130 4.280 ;
        RECT 502.970 0.155 505.350 4.280 ;
        RECT 506.190 0.155 508.570 4.280 ;
        RECT 509.410 0.155 511.790 4.280 ;
        RECT 512.630 0.155 515.010 4.280 ;
        RECT 515.850 0.155 518.230 4.280 ;
        RECT 519.070 0.155 521.450 4.280 ;
        RECT 522.290 0.155 524.670 4.280 ;
        RECT 525.510 0.155 527.890 4.280 ;
        RECT 528.730 0.155 531.110 4.280 ;
        RECT 531.950 0.155 534.330 4.280 ;
        RECT 535.170 0.155 537.550 4.280 ;
        RECT 538.390 0.155 540.770 4.280 ;
        RECT 541.610 0.155 543.990 4.280 ;
        RECT 544.830 0.155 547.210 4.280 ;
        RECT 548.050 0.155 550.430 4.280 ;
        RECT 551.270 0.155 553.650 4.280 ;
        RECT 554.490 0.155 556.870 4.280 ;
        RECT 557.710 0.155 560.090 4.280 ;
        RECT 560.930 0.155 563.310 4.280 ;
        RECT 564.150 0.155 566.530 4.280 ;
        RECT 567.370 0.155 569.750 4.280 ;
        RECT 570.590 0.155 572.970 4.280 ;
        RECT 573.810 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 582.630 4.280 ;
        RECT 583.470 0.155 585.850 4.280 ;
        RECT 586.690 0.155 589.070 4.280 ;
        RECT 589.910 0.155 592.290 4.280 ;
        RECT 593.130 0.155 595.510 4.280 ;
        RECT 596.350 0.155 598.730 4.280 ;
        RECT 599.570 0.155 601.950 4.280 ;
        RECT 602.790 0.155 605.170 4.280 ;
        RECT 606.010 0.155 608.390 4.280 ;
        RECT 609.230 0.155 611.610 4.280 ;
        RECT 612.450 0.155 614.830 4.280 ;
        RECT 615.670 0.155 618.050 4.280 ;
        RECT 618.890 0.155 621.270 4.280 ;
        RECT 622.110 0.155 624.490 4.280 ;
        RECT 625.330 0.155 627.710 4.280 ;
        RECT 628.550 0.155 630.930 4.280 ;
        RECT 631.770 0.155 634.150 4.280 ;
        RECT 634.990 0.155 637.370 4.280 ;
        RECT 638.210 0.155 640.590 4.280 ;
        RECT 641.430 0.155 643.810 4.280 ;
        RECT 644.650 0.155 647.030 4.280 ;
        RECT 647.870 0.155 650.250 4.280 ;
        RECT 651.090 0.155 653.470 4.280 ;
        RECT 654.310 0.155 656.690 4.280 ;
        RECT 657.530 0.155 659.910 4.280 ;
        RECT 660.750 0.155 663.130 4.280 ;
        RECT 663.970 0.155 666.350 4.280 ;
        RECT 667.190 0.155 669.570 4.280 ;
        RECT 670.410 0.155 672.790 4.280 ;
        RECT 673.630 0.155 676.010 4.280 ;
        RECT 676.850 0.155 679.230 4.280 ;
        RECT 680.070 0.155 682.450 4.280 ;
        RECT 683.290 0.155 685.670 4.280 ;
        RECT 686.510 0.155 688.890 4.280 ;
        RECT 689.730 0.155 692.110 4.280 ;
        RECT 692.950 0.155 695.330 4.280 ;
        RECT 696.170 0.155 698.550 4.280 ;
        RECT 699.390 0.155 701.770 4.280 ;
        RECT 702.610 0.155 704.990 4.280 ;
        RECT 705.830 0.155 708.210 4.280 ;
        RECT 709.050 0.155 711.430 4.280 ;
        RECT 712.270 0.155 714.650 4.280 ;
        RECT 715.490 0.155 717.870 4.280 ;
        RECT 718.710 0.155 721.090 4.280 ;
        RECT 721.930 0.155 724.310 4.280 ;
        RECT 725.150 0.155 727.530 4.280 ;
        RECT 728.370 0.155 730.750 4.280 ;
        RECT 731.590 0.155 733.970 4.280 ;
        RECT 734.810 0.155 737.190 4.280 ;
        RECT 738.030 0.155 740.410 4.280 ;
        RECT 741.250 0.155 743.630 4.280 ;
        RECT 744.470 0.155 746.850 4.280 ;
        RECT 747.690 0.155 750.070 4.280 ;
        RECT 750.910 0.155 753.290 4.280 ;
        RECT 754.130 0.155 756.510 4.280 ;
        RECT 757.350 0.155 759.730 4.280 ;
        RECT 760.570 0.155 762.950 4.280 ;
        RECT 763.790 0.155 766.170 4.280 ;
        RECT 767.010 0.155 769.390 4.280 ;
        RECT 770.230 0.155 772.610 4.280 ;
        RECT 773.450 0.155 775.830 4.280 ;
        RECT 776.670 0.155 779.050 4.280 ;
        RECT 779.890 0.155 782.270 4.280 ;
        RECT 783.110 0.155 785.490 4.280 ;
        RECT 786.330 0.155 788.710 4.280 ;
        RECT 789.550 0.155 791.930 4.280 ;
        RECT 792.770 0.155 795.150 4.280 ;
        RECT 795.990 0.155 798.370 4.280 ;
      LAYER met3 ;
        RECT 1.905 890.440 795.600 891.305 ;
        RECT 1.905 888.440 796.000 890.440 ;
        RECT 1.905 887.040 795.600 888.440 ;
        RECT 1.905 885.040 796.000 887.040 ;
        RECT 1.905 883.640 795.600 885.040 ;
        RECT 1.905 881.640 796.000 883.640 ;
        RECT 4.400 880.240 795.600 881.640 ;
        RECT 1.905 878.240 796.000 880.240 ;
        RECT 4.400 876.840 795.600 878.240 ;
        RECT 1.905 874.840 796.000 876.840 ;
        RECT 1.905 873.440 795.600 874.840 ;
        RECT 1.905 871.440 796.000 873.440 ;
        RECT 1.905 870.040 795.600 871.440 ;
        RECT 1.905 868.040 796.000 870.040 ;
        RECT 4.400 866.640 795.600 868.040 ;
        RECT 1.905 864.640 796.000 866.640 ;
        RECT 4.400 863.240 795.600 864.640 ;
        RECT 1.905 861.240 796.000 863.240 ;
        RECT 4.400 859.840 795.600 861.240 ;
        RECT 1.905 857.840 796.000 859.840 ;
        RECT 4.400 856.440 795.600 857.840 ;
        RECT 1.905 854.440 796.000 856.440 ;
        RECT 4.400 853.040 795.600 854.440 ;
        RECT 1.905 851.040 796.000 853.040 ;
        RECT 4.400 849.640 795.600 851.040 ;
        RECT 1.905 847.640 796.000 849.640 ;
        RECT 4.400 846.240 795.600 847.640 ;
        RECT 1.905 844.240 796.000 846.240 ;
        RECT 4.400 842.840 795.600 844.240 ;
        RECT 1.905 840.840 796.000 842.840 ;
        RECT 4.400 839.440 795.600 840.840 ;
        RECT 1.905 837.440 796.000 839.440 ;
        RECT 4.400 836.040 795.600 837.440 ;
        RECT 1.905 834.040 796.000 836.040 ;
        RECT 4.400 832.640 795.600 834.040 ;
        RECT 1.905 830.640 796.000 832.640 ;
        RECT 4.400 829.240 795.600 830.640 ;
        RECT 1.905 827.240 796.000 829.240 ;
        RECT 4.400 825.840 795.600 827.240 ;
        RECT 1.905 823.840 796.000 825.840 ;
        RECT 1.905 822.440 795.600 823.840 ;
        RECT 1.905 820.440 796.000 822.440 ;
        RECT 1.905 819.040 795.600 820.440 ;
        RECT 1.905 817.040 796.000 819.040 ;
        RECT 1.905 815.640 795.600 817.040 ;
        RECT 1.905 813.640 796.000 815.640 ;
        RECT 1.905 812.240 795.600 813.640 ;
        RECT 1.905 810.240 796.000 812.240 ;
        RECT 1.905 808.840 795.600 810.240 ;
        RECT 1.905 806.840 796.000 808.840 ;
        RECT 1.905 805.440 795.600 806.840 ;
        RECT 1.905 803.440 796.000 805.440 ;
        RECT 1.905 802.040 795.600 803.440 ;
        RECT 1.905 800.040 796.000 802.040 ;
        RECT 1.905 798.640 795.600 800.040 ;
        RECT 1.905 796.640 796.000 798.640 ;
        RECT 1.905 795.240 795.600 796.640 ;
        RECT 1.905 793.240 796.000 795.240 ;
        RECT 1.905 791.840 795.600 793.240 ;
        RECT 1.905 789.840 796.000 791.840 ;
        RECT 1.905 788.440 795.600 789.840 ;
        RECT 1.905 786.440 796.000 788.440 ;
        RECT 1.905 785.040 795.600 786.440 ;
        RECT 1.905 783.040 796.000 785.040 ;
        RECT 1.905 781.640 795.600 783.040 ;
        RECT 1.905 779.640 796.000 781.640 ;
        RECT 1.905 778.240 795.600 779.640 ;
        RECT 1.905 776.240 796.000 778.240 ;
        RECT 1.905 774.840 795.600 776.240 ;
        RECT 1.905 772.840 796.000 774.840 ;
        RECT 1.905 771.440 795.600 772.840 ;
        RECT 1.905 769.440 796.000 771.440 ;
        RECT 1.905 768.040 795.600 769.440 ;
        RECT 1.905 766.040 796.000 768.040 ;
        RECT 1.905 764.640 795.600 766.040 ;
        RECT 1.905 762.640 796.000 764.640 ;
        RECT 1.905 761.240 795.600 762.640 ;
        RECT 1.905 759.240 796.000 761.240 ;
        RECT 1.905 757.840 795.600 759.240 ;
        RECT 1.905 755.840 796.000 757.840 ;
        RECT 1.905 754.440 795.600 755.840 ;
        RECT 1.905 752.440 796.000 754.440 ;
        RECT 1.905 751.040 795.600 752.440 ;
        RECT 1.905 749.040 796.000 751.040 ;
        RECT 1.905 747.640 795.600 749.040 ;
        RECT 1.905 745.640 796.000 747.640 ;
        RECT 1.905 744.240 795.600 745.640 ;
        RECT 1.905 742.240 796.000 744.240 ;
        RECT 1.905 740.840 795.600 742.240 ;
        RECT 1.905 738.840 796.000 740.840 ;
        RECT 1.905 737.440 795.600 738.840 ;
        RECT 1.905 735.440 796.000 737.440 ;
        RECT 1.905 734.040 795.600 735.440 ;
        RECT 1.905 732.040 796.000 734.040 ;
        RECT 1.905 730.640 795.600 732.040 ;
        RECT 1.905 728.640 796.000 730.640 ;
        RECT 1.905 727.240 795.600 728.640 ;
        RECT 1.905 725.240 796.000 727.240 ;
        RECT 1.905 723.840 795.600 725.240 ;
        RECT 1.905 721.840 796.000 723.840 ;
        RECT 1.905 720.440 795.600 721.840 ;
        RECT 1.905 718.440 796.000 720.440 ;
        RECT 1.905 717.040 795.600 718.440 ;
        RECT 1.905 715.040 796.000 717.040 ;
        RECT 1.905 713.640 795.600 715.040 ;
        RECT 1.905 711.640 796.000 713.640 ;
        RECT 1.905 710.240 795.600 711.640 ;
        RECT 1.905 708.240 796.000 710.240 ;
        RECT 1.905 706.840 795.600 708.240 ;
        RECT 1.905 704.840 796.000 706.840 ;
        RECT 1.905 703.440 795.600 704.840 ;
        RECT 1.905 701.440 796.000 703.440 ;
        RECT 4.400 700.040 795.600 701.440 ;
        RECT 1.905 698.040 796.000 700.040 ;
        RECT 1.905 696.640 795.600 698.040 ;
        RECT 1.905 694.640 796.000 696.640 ;
        RECT 1.905 693.240 795.600 694.640 ;
        RECT 1.905 691.240 796.000 693.240 ;
        RECT 1.905 689.840 795.600 691.240 ;
        RECT 1.905 687.840 796.000 689.840 ;
        RECT 1.905 686.440 795.600 687.840 ;
        RECT 1.905 684.440 796.000 686.440 ;
        RECT 1.905 683.040 795.600 684.440 ;
        RECT 1.905 681.040 796.000 683.040 ;
        RECT 1.905 679.640 795.600 681.040 ;
        RECT 1.905 677.640 796.000 679.640 ;
        RECT 1.905 676.240 795.600 677.640 ;
        RECT 1.905 674.240 796.000 676.240 ;
        RECT 1.905 672.840 795.600 674.240 ;
        RECT 1.905 670.840 796.000 672.840 ;
        RECT 1.905 669.440 795.600 670.840 ;
        RECT 1.905 667.440 796.000 669.440 ;
        RECT 1.905 666.040 795.600 667.440 ;
        RECT 1.905 664.040 796.000 666.040 ;
        RECT 1.905 662.640 795.600 664.040 ;
        RECT 1.905 660.640 796.000 662.640 ;
        RECT 1.905 659.240 795.600 660.640 ;
        RECT 1.905 657.240 796.000 659.240 ;
        RECT 1.905 655.840 795.600 657.240 ;
        RECT 1.905 653.840 796.000 655.840 ;
        RECT 1.905 652.440 795.600 653.840 ;
        RECT 1.905 650.440 796.000 652.440 ;
        RECT 1.905 649.040 795.600 650.440 ;
        RECT 1.905 647.040 796.000 649.040 ;
        RECT 1.905 645.640 795.600 647.040 ;
        RECT 1.905 643.640 796.000 645.640 ;
        RECT 1.905 642.240 795.600 643.640 ;
        RECT 1.905 640.240 796.000 642.240 ;
        RECT 1.905 638.840 795.600 640.240 ;
        RECT 1.905 636.840 796.000 638.840 ;
        RECT 1.905 635.440 795.600 636.840 ;
        RECT 1.905 633.440 796.000 635.440 ;
        RECT 1.905 632.040 795.600 633.440 ;
        RECT 1.905 630.040 796.000 632.040 ;
        RECT 1.905 628.640 795.600 630.040 ;
        RECT 1.905 626.640 796.000 628.640 ;
        RECT 1.905 625.240 795.600 626.640 ;
        RECT 1.905 623.240 796.000 625.240 ;
        RECT 1.905 621.840 795.600 623.240 ;
        RECT 1.905 619.840 796.000 621.840 ;
        RECT 1.905 618.440 795.600 619.840 ;
        RECT 1.905 616.440 796.000 618.440 ;
        RECT 1.905 615.040 795.600 616.440 ;
        RECT 1.905 613.040 796.000 615.040 ;
        RECT 1.905 611.640 795.600 613.040 ;
        RECT 1.905 609.640 796.000 611.640 ;
        RECT 1.905 608.240 795.600 609.640 ;
        RECT 1.905 606.240 796.000 608.240 ;
        RECT 1.905 604.840 795.600 606.240 ;
        RECT 1.905 602.840 796.000 604.840 ;
        RECT 1.905 601.440 795.600 602.840 ;
        RECT 1.905 599.440 796.000 601.440 ;
        RECT 1.905 598.040 795.600 599.440 ;
        RECT 1.905 596.040 796.000 598.040 ;
        RECT 1.905 594.640 795.600 596.040 ;
        RECT 1.905 592.640 796.000 594.640 ;
        RECT 1.905 591.240 795.600 592.640 ;
        RECT 1.905 589.240 796.000 591.240 ;
        RECT 1.905 587.840 795.600 589.240 ;
        RECT 1.905 585.840 796.000 587.840 ;
        RECT 1.905 584.440 795.600 585.840 ;
        RECT 1.905 582.440 796.000 584.440 ;
        RECT 1.905 581.040 795.600 582.440 ;
        RECT 1.905 579.040 796.000 581.040 ;
        RECT 1.905 577.640 795.600 579.040 ;
        RECT 1.905 575.640 796.000 577.640 ;
        RECT 1.905 574.240 795.600 575.640 ;
        RECT 1.905 572.240 796.000 574.240 ;
        RECT 1.905 570.840 795.600 572.240 ;
        RECT 1.905 568.840 796.000 570.840 ;
        RECT 1.905 567.440 795.600 568.840 ;
        RECT 1.905 565.440 796.000 567.440 ;
        RECT 1.905 564.040 795.600 565.440 ;
        RECT 1.905 562.040 796.000 564.040 ;
        RECT 1.905 560.640 795.600 562.040 ;
        RECT 1.905 558.640 796.000 560.640 ;
        RECT 1.905 557.240 795.600 558.640 ;
        RECT 1.905 555.240 796.000 557.240 ;
        RECT 1.905 553.840 795.600 555.240 ;
        RECT 1.905 551.840 796.000 553.840 ;
        RECT 1.905 550.440 795.600 551.840 ;
        RECT 1.905 548.440 796.000 550.440 ;
        RECT 1.905 547.040 795.600 548.440 ;
        RECT 1.905 545.040 796.000 547.040 ;
        RECT 1.905 543.640 795.600 545.040 ;
        RECT 1.905 541.640 796.000 543.640 ;
        RECT 1.905 540.240 795.600 541.640 ;
        RECT 1.905 538.240 796.000 540.240 ;
        RECT 1.905 536.840 795.600 538.240 ;
        RECT 1.905 534.840 796.000 536.840 ;
        RECT 1.905 533.440 795.600 534.840 ;
        RECT 1.905 531.440 796.000 533.440 ;
        RECT 1.905 530.040 795.600 531.440 ;
        RECT 1.905 528.040 796.000 530.040 ;
        RECT 1.905 526.640 795.600 528.040 ;
        RECT 1.905 524.640 796.000 526.640 ;
        RECT 1.905 523.240 795.600 524.640 ;
        RECT 1.905 521.240 796.000 523.240 ;
        RECT 1.905 519.840 795.600 521.240 ;
        RECT 1.905 517.840 796.000 519.840 ;
        RECT 1.905 516.440 795.600 517.840 ;
        RECT 1.905 514.440 796.000 516.440 ;
        RECT 1.905 513.040 795.600 514.440 ;
        RECT 1.905 511.040 796.000 513.040 ;
        RECT 1.905 509.640 795.600 511.040 ;
        RECT 1.905 507.640 796.000 509.640 ;
        RECT 1.905 506.240 795.600 507.640 ;
        RECT 1.905 504.240 796.000 506.240 ;
        RECT 1.905 502.840 795.600 504.240 ;
        RECT 1.905 500.840 796.000 502.840 ;
        RECT 1.905 499.440 795.600 500.840 ;
        RECT 1.905 497.440 796.000 499.440 ;
        RECT 1.905 496.040 795.600 497.440 ;
        RECT 1.905 494.040 796.000 496.040 ;
        RECT 1.905 492.640 795.600 494.040 ;
        RECT 1.905 490.640 796.000 492.640 ;
        RECT 1.905 489.240 795.600 490.640 ;
        RECT 1.905 487.240 796.000 489.240 ;
        RECT 1.905 485.840 795.600 487.240 ;
        RECT 1.905 483.840 796.000 485.840 ;
        RECT 1.905 482.440 795.600 483.840 ;
        RECT 1.905 480.440 796.000 482.440 ;
        RECT 1.905 479.040 795.600 480.440 ;
        RECT 1.905 477.040 796.000 479.040 ;
        RECT 1.905 475.640 795.600 477.040 ;
        RECT 1.905 473.640 796.000 475.640 ;
        RECT 1.905 472.240 795.600 473.640 ;
        RECT 1.905 470.240 796.000 472.240 ;
        RECT 1.905 468.840 795.600 470.240 ;
        RECT 1.905 466.840 796.000 468.840 ;
        RECT 1.905 465.440 795.600 466.840 ;
        RECT 1.905 463.440 796.000 465.440 ;
        RECT 1.905 462.040 795.600 463.440 ;
        RECT 1.905 460.040 796.000 462.040 ;
        RECT 1.905 458.640 795.600 460.040 ;
        RECT 1.905 456.640 796.000 458.640 ;
        RECT 1.905 455.240 795.600 456.640 ;
        RECT 1.905 453.240 796.000 455.240 ;
        RECT 1.905 451.840 795.600 453.240 ;
        RECT 1.905 449.840 796.000 451.840 ;
        RECT 1.905 448.440 795.600 449.840 ;
        RECT 1.905 446.440 796.000 448.440 ;
        RECT 1.905 445.040 795.600 446.440 ;
        RECT 1.905 443.040 796.000 445.040 ;
        RECT 1.905 441.640 795.600 443.040 ;
        RECT 1.905 439.640 796.000 441.640 ;
        RECT 1.905 438.240 795.600 439.640 ;
        RECT 1.905 436.240 796.000 438.240 ;
        RECT 1.905 434.840 795.600 436.240 ;
        RECT 1.905 432.840 796.000 434.840 ;
        RECT 1.905 431.440 795.600 432.840 ;
        RECT 1.905 429.440 796.000 431.440 ;
        RECT 1.905 428.040 795.600 429.440 ;
        RECT 1.905 426.040 796.000 428.040 ;
        RECT 1.905 424.640 795.600 426.040 ;
        RECT 1.905 422.640 796.000 424.640 ;
        RECT 1.905 421.240 795.600 422.640 ;
        RECT 1.905 419.240 796.000 421.240 ;
        RECT 1.905 417.840 795.600 419.240 ;
        RECT 1.905 415.840 796.000 417.840 ;
        RECT 1.905 414.440 795.600 415.840 ;
        RECT 1.905 412.440 796.000 414.440 ;
        RECT 1.905 411.040 795.600 412.440 ;
        RECT 1.905 409.040 796.000 411.040 ;
        RECT 1.905 407.640 795.600 409.040 ;
        RECT 1.905 405.640 796.000 407.640 ;
        RECT 1.905 404.240 795.600 405.640 ;
        RECT 1.905 402.240 796.000 404.240 ;
        RECT 1.905 400.840 795.600 402.240 ;
        RECT 1.905 398.840 796.000 400.840 ;
        RECT 1.905 397.440 795.600 398.840 ;
        RECT 1.905 395.440 796.000 397.440 ;
        RECT 1.905 394.040 795.600 395.440 ;
        RECT 1.905 392.040 796.000 394.040 ;
        RECT 1.905 390.640 795.600 392.040 ;
        RECT 1.905 388.640 796.000 390.640 ;
        RECT 1.905 387.240 795.600 388.640 ;
        RECT 1.905 385.240 796.000 387.240 ;
        RECT 1.905 383.840 795.600 385.240 ;
        RECT 1.905 381.840 796.000 383.840 ;
        RECT 1.905 380.440 795.600 381.840 ;
        RECT 1.905 378.440 796.000 380.440 ;
        RECT 1.905 377.040 795.600 378.440 ;
        RECT 1.905 375.040 796.000 377.040 ;
        RECT 1.905 373.640 795.600 375.040 ;
        RECT 1.905 371.640 796.000 373.640 ;
        RECT 1.905 370.240 795.600 371.640 ;
        RECT 1.905 368.240 796.000 370.240 ;
        RECT 1.905 366.840 795.600 368.240 ;
        RECT 1.905 364.840 796.000 366.840 ;
        RECT 1.905 363.440 795.600 364.840 ;
        RECT 1.905 361.440 796.000 363.440 ;
        RECT 1.905 360.040 795.600 361.440 ;
        RECT 1.905 358.040 796.000 360.040 ;
        RECT 1.905 356.640 795.600 358.040 ;
        RECT 1.905 354.640 796.000 356.640 ;
        RECT 1.905 353.240 795.600 354.640 ;
        RECT 1.905 351.240 796.000 353.240 ;
        RECT 1.905 349.840 795.600 351.240 ;
        RECT 1.905 347.840 796.000 349.840 ;
        RECT 1.905 346.440 795.600 347.840 ;
        RECT 1.905 344.440 796.000 346.440 ;
        RECT 1.905 343.040 795.600 344.440 ;
        RECT 1.905 341.040 796.000 343.040 ;
        RECT 1.905 339.640 795.600 341.040 ;
        RECT 1.905 337.640 796.000 339.640 ;
        RECT 1.905 336.240 795.600 337.640 ;
        RECT 1.905 334.240 796.000 336.240 ;
        RECT 1.905 332.840 795.600 334.240 ;
        RECT 1.905 330.840 796.000 332.840 ;
        RECT 1.905 329.440 795.600 330.840 ;
        RECT 1.905 327.440 796.000 329.440 ;
        RECT 1.905 326.040 795.600 327.440 ;
        RECT 1.905 324.040 796.000 326.040 ;
        RECT 1.905 322.640 795.600 324.040 ;
        RECT 1.905 320.640 796.000 322.640 ;
        RECT 1.905 319.240 795.600 320.640 ;
        RECT 1.905 317.240 796.000 319.240 ;
        RECT 1.905 315.840 795.600 317.240 ;
        RECT 1.905 313.840 796.000 315.840 ;
        RECT 1.905 312.440 795.600 313.840 ;
        RECT 1.905 310.440 796.000 312.440 ;
        RECT 1.905 309.040 795.600 310.440 ;
        RECT 1.905 307.040 796.000 309.040 ;
        RECT 1.905 305.640 795.600 307.040 ;
        RECT 1.905 303.640 796.000 305.640 ;
        RECT 1.905 302.240 795.600 303.640 ;
        RECT 1.905 300.240 796.000 302.240 ;
        RECT 1.905 298.840 795.600 300.240 ;
        RECT 1.905 296.840 796.000 298.840 ;
        RECT 1.905 295.440 795.600 296.840 ;
        RECT 1.905 293.440 796.000 295.440 ;
        RECT 1.905 292.040 795.600 293.440 ;
        RECT 1.905 290.040 796.000 292.040 ;
        RECT 1.905 288.640 795.600 290.040 ;
        RECT 1.905 286.640 796.000 288.640 ;
        RECT 1.905 285.240 795.600 286.640 ;
        RECT 1.905 283.240 796.000 285.240 ;
        RECT 1.905 281.840 795.600 283.240 ;
        RECT 1.905 279.840 796.000 281.840 ;
        RECT 1.905 278.440 795.600 279.840 ;
        RECT 1.905 276.440 796.000 278.440 ;
        RECT 1.905 275.040 795.600 276.440 ;
        RECT 1.905 273.040 796.000 275.040 ;
        RECT 1.905 271.640 795.600 273.040 ;
        RECT 1.905 269.640 796.000 271.640 ;
        RECT 1.905 268.240 795.600 269.640 ;
        RECT 1.905 266.240 796.000 268.240 ;
        RECT 1.905 264.840 795.600 266.240 ;
        RECT 1.905 262.840 796.000 264.840 ;
        RECT 1.905 261.440 795.600 262.840 ;
        RECT 1.905 259.440 796.000 261.440 ;
        RECT 1.905 258.040 795.600 259.440 ;
        RECT 1.905 256.040 796.000 258.040 ;
        RECT 1.905 254.640 795.600 256.040 ;
        RECT 1.905 252.640 796.000 254.640 ;
        RECT 1.905 251.240 795.600 252.640 ;
        RECT 1.905 249.240 796.000 251.240 ;
        RECT 1.905 247.840 795.600 249.240 ;
        RECT 1.905 245.840 796.000 247.840 ;
        RECT 1.905 244.440 795.600 245.840 ;
        RECT 1.905 242.440 796.000 244.440 ;
        RECT 1.905 241.040 795.600 242.440 ;
        RECT 1.905 239.040 796.000 241.040 ;
        RECT 1.905 237.640 795.600 239.040 ;
        RECT 1.905 235.640 796.000 237.640 ;
        RECT 1.905 234.240 795.600 235.640 ;
        RECT 1.905 232.240 796.000 234.240 ;
        RECT 1.905 230.840 795.600 232.240 ;
        RECT 1.905 228.840 796.000 230.840 ;
        RECT 1.905 227.440 795.600 228.840 ;
        RECT 1.905 225.440 796.000 227.440 ;
        RECT 1.905 224.040 795.600 225.440 ;
        RECT 1.905 222.040 796.000 224.040 ;
        RECT 1.905 220.640 795.600 222.040 ;
        RECT 1.905 218.640 796.000 220.640 ;
        RECT 1.905 217.240 795.600 218.640 ;
        RECT 1.905 215.240 796.000 217.240 ;
        RECT 1.905 213.840 795.600 215.240 ;
        RECT 1.905 211.840 796.000 213.840 ;
        RECT 1.905 210.440 795.600 211.840 ;
        RECT 1.905 208.440 796.000 210.440 ;
        RECT 1.905 207.040 795.600 208.440 ;
        RECT 1.905 205.040 796.000 207.040 ;
        RECT 1.905 203.640 795.600 205.040 ;
        RECT 1.905 201.640 796.000 203.640 ;
        RECT 1.905 200.240 795.600 201.640 ;
        RECT 1.905 198.240 796.000 200.240 ;
        RECT 1.905 196.840 795.600 198.240 ;
        RECT 1.905 194.840 796.000 196.840 ;
        RECT 1.905 193.440 795.600 194.840 ;
        RECT 1.905 191.440 796.000 193.440 ;
        RECT 1.905 190.040 795.600 191.440 ;
        RECT 1.905 188.040 796.000 190.040 ;
        RECT 1.905 186.640 795.600 188.040 ;
        RECT 1.905 184.640 796.000 186.640 ;
        RECT 1.905 183.240 795.600 184.640 ;
        RECT 1.905 181.240 796.000 183.240 ;
        RECT 1.905 179.840 795.600 181.240 ;
        RECT 1.905 177.840 796.000 179.840 ;
        RECT 1.905 176.440 795.600 177.840 ;
        RECT 1.905 174.440 796.000 176.440 ;
        RECT 1.905 173.040 795.600 174.440 ;
        RECT 1.905 171.040 796.000 173.040 ;
        RECT 1.905 169.640 795.600 171.040 ;
        RECT 1.905 167.640 796.000 169.640 ;
        RECT 1.905 166.240 795.600 167.640 ;
        RECT 1.905 164.240 796.000 166.240 ;
        RECT 1.905 162.840 795.600 164.240 ;
        RECT 1.905 160.840 796.000 162.840 ;
        RECT 1.905 159.440 795.600 160.840 ;
        RECT 1.905 157.440 796.000 159.440 ;
        RECT 1.905 156.040 795.600 157.440 ;
        RECT 1.905 154.040 796.000 156.040 ;
        RECT 1.905 152.640 795.600 154.040 ;
        RECT 1.905 150.640 796.000 152.640 ;
        RECT 1.905 149.240 795.600 150.640 ;
        RECT 1.905 147.240 796.000 149.240 ;
        RECT 1.905 145.840 795.600 147.240 ;
        RECT 1.905 143.840 796.000 145.840 ;
        RECT 1.905 142.440 795.600 143.840 ;
        RECT 1.905 140.440 796.000 142.440 ;
        RECT 1.905 139.040 795.600 140.440 ;
        RECT 1.905 137.040 796.000 139.040 ;
        RECT 4.400 135.640 795.600 137.040 ;
        RECT 1.905 133.640 796.000 135.640 ;
        RECT 1.905 132.240 795.600 133.640 ;
        RECT 1.905 130.240 796.000 132.240 ;
        RECT 1.905 128.840 795.600 130.240 ;
        RECT 1.905 126.840 796.000 128.840 ;
        RECT 1.905 125.440 795.600 126.840 ;
        RECT 1.905 123.440 796.000 125.440 ;
        RECT 1.905 122.040 795.600 123.440 ;
        RECT 1.905 120.040 796.000 122.040 ;
        RECT 1.905 118.640 795.600 120.040 ;
        RECT 1.905 116.640 796.000 118.640 ;
        RECT 1.905 115.240 795.600 116.640 ;
        RECT 1.905 113.240 796.000 115.240 ;
        RECT 1.905 111.840 795.600 113.240 ;
        RECT 1.905 109.840 796.000 111.840 ;
        RECT 4.400 108.440 795.600 109.840 ;
        RECT 1.905 106.440 796.000 108.440 ;
        RECT 1.905 105.040 795.600 106.440 ;
        RECT 1.905 103.040 796.000 105.040 ;
        RECT 1.905 101.640 795.600 103.040 ;
        RECT 1.905 99.640 796.000 101.640 ;
        RECT 1.905 98.240 795.600 99.640 ;
        RECT 1.905 96.240 796.000 98.240 ;
        RECT 1.905 94.840 795.600 96.240 ;
        RECT 1.905 92.840 796.000 94.840 ;
        RECT 1.905 91.440 795.600 92.840 ;
        RECT 1.905 89.440 796.000 91.440 ;
        RECT 1.905 88.040 795.600 89.440 ;
        RECT 1.905 86.040 796.000 88.040 ;
        RECT 1.905 84.640 795.600 86.040 ;
        RECT 1.905 82.640 796.000 84.640 ;
        RECT 1.905 81.240 795.600 82.640 ;
        RECT 1.905 79.240 796.000 81.240 ;
        RECT 1.905 77.840 795.600 79.240 ;
        RECT 1.905 75.840 796.000 77.840 ;
        RECT 1.905 74.440 795.600 75.840 ;
        RECT 1.905 72.440 796.000 74.440 ;
        RECT 1.905 71.040 795.600 72.440 ;
        RECT 1.905 69.040 796.000 71.040 ;
        RECT 4.400 67.640 795.600 69.040 ;
        RECT 1.905 65.640 796.000 67.640 ;
        RECT 1.905 64.240 795.600 65.640 ;
        RECT 1.905 62.240 796.000 64.240 ;
        RECT 1.905 60.840 795.600 62.240 ;
        RECT 1.905 58.840 796.000 60.840 ;
        RECT 1.905 57.440 795.600 58.840 ;
        RECT 1.905 55.440 796.000 57.440 ;
        RECT 4.400 54.040 795.600 55.440 ;
        RECT 1.905 52.040 796.000 54.040 ;
        RECT 1.905 50.640 795.600 52.040 ;
        RECT 1.905 48.640 796.000 50.640 ;
        RECT 1.905 47.240 795.600 48.640 ;
        RECT 1.905 45.240 796.000 47.240 ;
        RECT 4.400 43.840 795.600 45.240 ;
        RECT 1.905 41.840 796.000 43.840 ;
        RECT 4.400 40.440 795.600 41.840 ;
        RECT 1.905 38.440 796.000 40.440 ;
        RECT 1.905 37.040 795.600 38.440 ;
        RECT 1.905 35.040 796.000 37.040 ;
        RECT 1.905 33.640 795.600 35.040 ;
        RECT 1.905 31.640 796.000 33.640 ;
        RECT 1.905 30.240 795.600 31.640 ;
        RECT 1.905 28.240 796.000 30.240 ;
        RECT 1.905 26.840 795.600 28.240 ;
        RECT 1.905 24.840 796.000 26.840 ;
        RECT 4.400 23.440 795.600 24.840 ;
        RECT 1.905 21.440 796.000 23.440 ;
        RECT 1.905 20.040 795.600 21.440 ;
        RECT 1.905 18.040 796.000 20.040 ;
        RECT 4.400 16.640 795.600 18.040 ;
        RECT 1.905 14.640 796.000 16.640 ;
        RECT 1.905 13.240 795.600 14.640 ;
        RECT 1.905 11.240 796.000 13.240 ;
        RECT 1.905 9.840 795.600 11.240 ;
        RECT 1.905 7.840 796.000 9.840 ;
        RECT 1.905 6.440 795.600 7.840 ;
        RECT 1.905 4.440 796.000 6.440 ;
        RECT 1.905 3.040 795.600 4.440 ;
        RECT 1.905 1.040 796.000 3.040 ;
        RECT 1.905 0.175 795.600 1.040 ;
      LAYER met4 ;
        RECT 5.815 17.175 20.640 885.865 ;
        RECT 23.040 17.175 23.940 885.865 ;
        RECT 26.340 17.175 174.240 885.865 ;
        RECT 176.640 17.175 177.540 885.865 ;
        RECT 179.940 17.175 327.840 885.865 ;
        RECT 330.240 17.175 331.140 885.865 ;
        RECT 333.540 17.175 481.440 885.865 ;
        RECT 483.840 17.175 484.740 885.865 ;
        RECT 487.140 17.175 635.040 885.865 ;
        RECT 637.440 17.175 638.340 885.865 ;
        RECT 640.740 17.175 786.305 885.865 ;
  END
END team_12_Wrapper
END LIBRARY

