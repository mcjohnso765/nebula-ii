VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO team_03
  CLASS BLOCK ;
  FOREIGN team_03 ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 400.000 ;
  PIN ACK_I
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.970 396.000 13.250 400.000 ;
    END
  END ACK_I
  PIN ADR_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 396.000 267.630 400.000 ;
    END
  END ADR_O[0]
  PIN ADR_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 389.710 396.000 389.990 400.000 ;
    END
  END ADR_O[10]
  PIN ADR_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 396.150 396.000 396.430 400.000 ;
    END
  END ADR_O[11]
  PIN ADR_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 412.250 396.000 412.530 400.000 ;
    END
  END ADR_O[12]
  PIN ADR_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 447.670 396.000 447.950 400.000 ;
    END
  END ADR_O[13]
  PIN ADR_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 431.570 396.000 431.850 400.000 ;
    END
  END ADR_O[14]
  PIN ADR_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 470.210 396.000 470.490 400.000 ;
    END
  END ADR_O[15]
  PIN ADR_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 486.310 396.000 486.590 400.000 ;
    END
  END ADR_O[16]
  PIN ADR_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 502.410 396.000 502.690 400.000 ;
    END
  END ADR_O[17]
  PIN ADR_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 396.000 325.590 400.000 ;
    END
  END ADR_O[18]
  PIN ADR_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 396.000 335.250 400.000 ;
    END
  END ADR_O[19]
  PIN ADR_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 396.000 254.750 400.000 ;
    END
  END ADR_O[1]
  PIN ADR_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 396.000 312.710 400.000 ;
    END
  END ADR_O[20]
  PIN ADR_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 396.000 299.830 400.000 ;
    END
  END ADR_O[21]
  PIN ADR_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 283.450 396.000 283.730 400.000 ;
    END
  END ADR_O[22]
  PIN ADR_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 270.570 396.000 270.850 400.000 ;
    END
  END ADR_O[23]
  PIN ADR_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 396.000 241.870 400.000 ;
    END
  END ADR_O[24]
  PIN ADR_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 396.000 225.770 400.000 ;
    END
  END ADR_O[25]
  PIN ADR_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 396.000 219.330 400.000 ;
    END
  END ADR_O[26]
  PIN ADR_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.310 396.000 3.590 400.000 ;
    END
  END ADR_O[27]
  PIN ADR_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 396.000 42.230 400.000 ;
    END
  END ADR_O[28]
  PIN ADR_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 396.000 48.670 400.000 ;
    END
  END ADR_O[29]
  PIN ADR_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 570.030 396.000 570.310 400.000 ;
    END
  END ADR_O[2]
  PIN ADR_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 396.000 6.810 400.000 ;
    END
  END ADR_O[30]
  PIN ADR_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 396.000 10.030 400.000 ;
    END
  END ADR_O[31]
  PIN ADR_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 560.370 396.000 560.650 400.000 ;
    END
  END ADR_O[3]
  PIN ADR_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 541.050 396.000 541.330 400.000 ;
    END
  END ADR_O[4]
  PIN ADR_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 563.590 396.000 563.870 400.000 ;
    END
  END ADR_O[5]
  PIN ADR_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 524.950 396.000 525.230 400.000 ;
    END
  END ADR_O[6]
  PIN ADR_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 515.290 396.000 515.570 400.000 ;
    END
  END ADR_O[7]
  PIN ADR_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 396.000 370.670 400.000 ;
    END
  END ADR_O[8]
  PIN ADR_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 354.290 396.000 354.570 400.000 ;
    END
  END ADR_O[9]
  PIN CYC_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 396.000 16.470 400.000 ;
    END
  END CYC_O
  PIN DAT_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 396.000 39.010 400.000 ;
    END
  END DAT_I[0]
  PIN DAT_I[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END DAT_I[10]
  PIN DAT_I[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END DAT_I[11]
  PIN DAT_I[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END DAT_I[12]
  PIN DAT_I[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 396.000 19.690 400.000 ;
    END
  END DAT_I[13]
  PIN DAT_I[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END DAT_I[14]
  PIN DAT_I[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END DAT_I[15]
  PIN DAT_I[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END DAT_I[16]
  PIN DAT_I[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.510 396.000 35.790 400.000 ;
    END
  END DAT_I[17]
  PIN DAT_I[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END DAT_I[18]
  PIN DAT_I[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END DAT_I[19]
  PIN DAT_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 396.000 32.570 400.000 ;
    END
  END DAT_I[1]
  PIN DAT_I[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END DAT_I[20]
  PIN DAT_I[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END DAT_I[21]
  PIN DAT_I[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END DAT_I[22]
  PIN DAT_I[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 0.090 396.000 0.370 400.000 ;
    END
  END DAT_I[23]
  PIN DAT_I[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END DAT_I[24]
  PIN DAT_I[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 396.000 45.450 400.000 ;
    END
  END DAT_I[25]
  PIN DAT_I[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.630 396.000 22.910 400.000 ;
    END
  END DAT_I[26]
  PIN DAT_I[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 396.000 29.350 400.000 ;
    END
  END DAT_I[27]
  PIN DAT_I[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.830 396.000 55.110 400.000 ;
    END
  END DAT_I[28]
  PIN DAT_I[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 396.000 51.890 400.000 ;
    END
  END DAT_I[29]
  PIN DAT_I[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END DAT_I[2]
  PIN DAT_I[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 25.850 396.000 26.130 400.000 ;
    END
  END DAT_I[30]
  PIN DAT_I[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END DAT_I[31]
  PIN DAT_I[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END DAT_I[3]
  PIN DAT_I[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END DAT_I[4]
  PIN DAT_I[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END DAT_I[5]
  PIN DAT_I[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END DAT_I[6]
  PIN DAT_I[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END DAT_I[7]
  PIN DAT_I[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END DAT_I[8]
  PIN DAT_I[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END DAT_I[9]
  PIN DAT_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 696.000 397.840 700.000 398.440 ;
    END
  END DAT_O[0]
  PIN DAT_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 95.240 700.000 95.840 ;
    END
  END DAT_O[10]
  PIN DAT_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 105.440 700.000 106.040 ;
    END
  END DAT_O[11]
  PIN DAT_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 112.240 700.000 112.840 ;
    END
  END DAT_O[12]
  PIN DAT_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 180.240 700.000 180.840 ;
    END
  END DAT_O[13]
  PIN DAT_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 146.240 700.000 146.840 ;
    END
  END DAT_O[14]
  PIN DAT_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 149.640 700.000 150.240 ;
    END
  END DAT_O[15]
  PIN DAT_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 200.640 700.000 201.240 ;
    END
  END DAT_O[16]
  PIN DAT_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 265.240 700.000 265.840 ;
    END
  END DAT_O[17]
  PIN DAT_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 370.640 700.000 371.240 ;
    END
  END DAT_O[18]
  PIN DAT_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 98.640 700.000 99.240 ;
    END
  END DAT_O[19]
  PIN DAT_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 119.040 700.000 119.640 ;
    END
  END DAT_O[1]
  PIN DAT_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 217.640 700.000 218.240 ;
    END
  END DAT_O[20]
  PIN DAT_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 272.040 700.000 272.640 ;
    END
  END DAT_O[21]
  PIN DAT_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 268.640 700.000 269.240 ;
    END
  END DAT_O[22]
  PIN DAT_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 380.840 700.000 381.440 ;
    END
  END DAT_O[23]
  PIN DAT_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 329.840 700.000 330.440 ;
    END
  END DAT_O[24]
  PIN DAT_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 323.040 700.000 323.640 ;
    END
  END DAT_O[25]
  PIN DAT_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 261.840 700.000 262.440 ;
    END
  END DAT_O[26]
  PIN DAT_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 479.870 396.000 480.150 400.000 ;
    END
  END DAT_O[27]
  PIN DAT_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 326.440 700.000 327.040 ;
    END
  END DAT_O[28]
  PIN DAT_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 360.440 700.000 361.040 ;
    END
  END DAT_O[29]
  PIN DAT_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 166.640 700.000 167.240 ;
    END
  END DAT_O[2]
  PIN DAT_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 391.040 700.000 391.640 ;
    END
  END DAT_O[30]
  PIN DAT_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 224.440 700.000 225.040 ;
    END
  END DAT_O[31]
  PIN DAT_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 153.040 700.000 153.640 ;
    END
  END DAT_O[3]
  PIN DAT_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 163.240 700.000 163.840 ;
    END
  END DAT_O[4]
  PIN DAT_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 142.840 700.000 143.440 ;
    END
  END DAT_O[5]
  PIN DAT_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 136.040 700.000 136.640 ;
    END
  END DAT_O[6]
  PIN DAT_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 214.240 700.000 214.840 ;
    END
  END DAT_O[7]
  PIN DAT_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 132.640 700.000 133.240 ;
    END
  END DAT_O[8]
  PIN DAT_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 374.040 700.000 374.640 ;
    END
  END DAT_O[9]
  PIN SEL_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 396.000 145.270 400.000 ;
    END
  END SEL_O[0]
  PIN SEL_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 396.000 138.830 400.000 ;
    END
  END SEL_O[1]
  PIN SEL_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 396.000 142.050 400.000 ;
    END
  END SEL_O[2]
  PIN SEL_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 396.000 135.610 400.000 ;
    END
  END SEL_O[3]
  PIN STB_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END STB_O
  PIN WE_O
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 353.640 700.000 354.240 ;
    END
  END WE_O
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END en
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 289.890 396.000 290.170 400.000 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 257.690 396.000 257.970 400.000 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 396.000 296.610 400.000 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 273.790 396.000 274.070 400.000 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 396.000 338.470 400.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 331.750 396.000 332.030 400.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.130 396.000 264.410 400.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 277.010 396.000 277.290 400.000 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END gpio_in[33]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 260.910 396.000 261.190 400.000 ;
    END
  END gpio_in[3]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 302.770 396.000 303.050 400.000 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 286.670 396.000 286.950 400.000 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END gpio_in[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 336.640 700.000 337.240 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 231.240 700.000 231.840 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 125.840 700.000 126.440 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 122.440 700.000 123.040 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 176.840 700.000 177.440 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 278.840 700.000 279.440 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 159.840 700.000 160.440 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 183.640 700.000 184.240 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 207.440 700.000 208.040 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 367.240 700.000 367.840 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 302.640 700.000 303.240 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 299.240 700.000 299.840 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 495.970 396.000 496.250 400.000 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 258.440 700.000 259.040 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 492.750 396.000 493.030 400.000 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 387.640 700.000 388.240 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 333.240 700.000 333.840 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 319.640 700.000 320.240 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 197.240 700.000 197.840 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 460.550 396.000 460.830 400.000 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 312.840 700.000 313.440 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 696.000 394.440 700.000 395.040 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 241.440 700.000 242.040 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 102.040 700.000 102.640 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 244.840 700.000 245.440 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 275.440 700.000 276.040 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 238.040 700.000 238.640 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 255.040 700.000 255.640 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 285.640 700.000 286.240 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 251.640 700.000 252.240 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 129.240 700.000 129.840 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 343.440 700.000 344.040 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 309.440 700.000 310.040 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 234.640 700.000 235.240 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.840 700.000 296.440 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 115.640 700.000 116.240 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 173.440 700.000 174.040 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 282.240 700.000 282.840 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 156.440 700.000 157.040 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 187.040 700.000 187.640 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 193.840 700.000 194.440 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 363.840 700.000 364.440 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 306.040 700.000 306.640 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 108.840 700.000 109.440 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 489.530 396.000 489.810 400.000 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 204.040 700.000 204.640 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 505.630 396.000 505.910 400.000 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 384.240 700.000 384.840 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 340.040 700.000 340.640 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 316.240 700.000 316.840 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 190.440 700.000 191.040 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 457.330 396.000 457.610 400.000 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 346.840 700.000 347.440 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 350.240 700.000 350.840 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 221.040 700.000 221.640 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 357.040 700.000 357.640 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 248.240 700.000 248.840 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END gpio_out[33]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 170.040 700.000 170.640 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 210.840 700.000 211.440 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 289.040 700.000 289.640 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 139.440 700.000 140.040 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 227.840 700.000 228.440 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 292.440 700.000 293.040 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 377.440 700.000 378.040 ;
    END
  END gpio_out[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 34.040 700.000 34.640 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 389.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 694.330 389.150 ;
      LAYER li1 ;
        RECT 5.520 10.795 694.140 389.045 ;
      LAYER met1 ;
        RECT 0.070 10.640 694.440 390.280 ;
      LAYER met2 ;
        RECT 0.650 395.720 3.030 398.325 ;
        RECT 3.870 395.720 6.250 398.325 ;
        RECT 7.090 395.720 9.470 398.325 ;
        RECT 10.310 395.720 12.690 398.325 ;
        RECT 13.530 395.720 15.910 398.325 ;
        RECT 16.750 395.720 19.130 398.325 ;
        RECT 19.970 395.720 22.350 398.325 ;
        RECT 23.190 395.720 25.570 398.325 ;
        RECT 26.410 395.720 28.790 398.325 ;
        RECT 29.630 395.720 32.010 398.325 ;
        RECT 32.850 395.720 35.230 398.325 ;
        RECT 36.070 395.720 38.450 398.325 ;
        RECT 39.290 395.720 41.670 398.325 ;
        RECT 42.510 395.720 44.890 398.325 ;
        RECT 45.730 395.720 48.110 398.325 ;
        RECT 48.950 395.720 51.330 398.325 ;
        RECT 52.170 395.720 54.550 398.325 ;
        RECT 55.390 395.720 135.050 398.325 ;
        RECT 135.890 395.720 138.270 398.325 ;
        RECT 139.110 395.720 141.490 398.325 ;
        RECT 142.330 395.720 144.710 398.325 ;
        RECT 145.550 395.720 218.770 398.325 ;
        RECT 219.610 395.720 225.210 398.325 ;
        RECT 226.050 395.720 241.310 398.325 ;
        RECT 242.150 395.720 254.190 398.325 ;
        RECT 255.030 395.720 257.410 398.325 ;
        RECT 258.250 395.720 260.630 398.325 ;
        RECT 261.470 395.720 263.850 398.325 ;
        RECT 264.690 395.720 267.070 398.325 ;
        RECT 267.910 395.720 270.290 398.325 ;
        RECT 271.130 395.720 273.510 398.325 ;
        RECT 274.350 395.720 276.730 398.325 ;
        RECT 277.570 395.720 283.170 398.325 ;
        RECT 284.010 395.720 286.390 398.325 ;
        RECT 287.230 395.720 289.610 398.325 ;
        RECT 290.450 395.720 296.050 398.325 ;
        RECT 296.890 395.720 299.270 398.325 ;
        RECT 300.110 395.720 302.490 398.325 ;
        RECT 303.330 395.720 312.150 398.325 ;
        RECT 312.990 395.720 325.030 398.325 ;
        RECT 325.870 395.720 331.470 398.325 ;
        RECT 332.310 395.720 334.690 398.325 ;
        RECT 335.530 395.720 337.910 398.325 ;
        RECT 338.750 395.720 354.010 398.325 ;
        RECT 354.850 395.720 370.110 398.325 ;
        RECT 370.950 395.720 389.430 398.325 ;
        RECT 390.270 395.720 395.870 398.325 ;
        RECT 396.710 395.720 411.970 398.325 ;
        RECT 412.810 395.720 431.290 398.325 ;
        RECT 432.130 395.720 447.390 398.325 ;
        RECT 448.230 395.720 457.050 398.325 ;
        RECT 457.890 395.720 460.270 398.325 ;
        RECT 461.110 395.720 469.930 398.325 ;
        RECT 470.770 395.720 479.590 398.325 ;
        RECT 480.430 395.720 486.030 398.325 ;
        RECT 486.870 395.720 489.250 398.325 ;
        RECT 490.090 395.720 492.470 398.325 ;
        RECT 493.310 395.720 495.690 398.325 ;
        RECT 496.530 395.720 502.130 398.325 ;
        RECT 502.970 395.720 505.350 398.325 ;
        RECT 506.190 395.720 515.010 398.325 ;
        RECT 515.850 395.720 524.670 398.325 ;
        RECT 525.510 395.720 540.770 398.325 ;
        RECT 541.610 395.720 560.090 398.325 ;
        RECT 560.930 395.720 563.310 398.325 ;
        RECT 564.150 395.720 569.750 398.325 ;
        RECT 570.590 395.720 693.590 398.325 ;
        RECT 0.100 10.695 693.590 395.720 ;
      LAYER met3 ;
        RECT 3.990 397.440 695.600 398.305 ;
        RECT 3.990 395.440 696.000 397.440 ;
        RECT 3.990 394.040 695.600 395.440 ;
        RECT 3.990 392.040 696.000 394.040 ;
        RECT 3.990 390.640 695.600 392.040 ;
        RECT 3.990 388.640 696.000 390.640 ;
        RECT 3.990 387.240 695.600 388.640 ;
        RECT 3.990 385.240 696.000 387.240 ;
        RECT 3.990 383.840 695.600 385.240 ;
        RECT 3.990 381.840 696.000 383.840 ;
        RECT 4.400 380.440 695.600 381.840 ;
        RECT 3.990 378.440 696.000 380.440 ;
        RECT 4.400 377.040 695.600 378.440 ;
        RECT 3.990 375.040 696.000 377.040 ;
        RECT 4.400 373.640 695.600 375.040 ;
        RECT 3.990 371.640 696.000 373.640 ;
        RECT 4.400 370.240 695.600 371.640 ;
        RECT 3.990 368.240 696.000 370.240 ;
        RECT 4.400 366.840 695.600 368.240 ;
        RECT 3.990 364.840 696.000 366.840 ;
        RECT 4.400 363.440 695.600 364.840 ;
        RECT 3.990 361.440 696.000 363.440 ;
        RECT 4.400 360.040 695.600 361.440 ;
        RECT 3.990 358.040 696.000 360.040 ;
        RECT 3.990 356.640 695.600 358.040 ;
        RECT 3.990 354.640 696.000 356.640 ;
        RECT 3.990 353.240 695.600 354.640 ;
        RECT 3.990 351.240 696.000 353.240 ;
        RECT 4.400 349.840 695.600 351.240 ;
        RECT 3.990 347.840 696.000 349.840 ;
        RECT 4.400 346.440 695.600 347.840 ;
        RECT 3.990 344.440 696.000 346.440 ;
        RECT 4.400 343.040 695.600 344.440 ;
        RECT 3.990 341.040 696.000 343.040 ;
        RECT 4.400 339.640 695.600 341.040 ;
        RECT 3.990 337.640 696.000 339.640 ;
        RECT 4.400 336.240 695.600 337.640 ;
        RECT 3.990 334.240 696.000 336.240 ;
        RECT 4.400 332.840 695.600 334.240 ;
        RECT 3.990 330.840 696.000 332.840 ;
        RECT 4.400 329.440 695.600 330.840 ;
        RECT 3.990 327.440 696.000 329.440 ;
        RECT 4.400 326.040 695.600 327.440 ;
        RECT 3.990 324.040 696.000 326.040 ;
        RECT 4.400 322.640 695.600 324.040 ;
        RECT 3.990 320.640 696.000 322.640 ;
        RECT 4.400 319.240 695.600 320.640 ;
        RECT 3.990 317.240 696.000 319.240 ;
        RECT 4.400 315.840 695.600 317.240 ;
        RECT 3.990 313.840 696.000 315.840 ;
        RECT 4.400 312.440 695.600 313.840 ;
        RECT 3.990 310.440 696.000 312.440 ;
        RECT 4.400 309.040 695.600 310.440 ;
        RECT 3.990 307.040 696.000 309.040 ;
        RECT 4.400 305.640 695.600 307.040 ;
        RECT 3.990 303.640 696.000 305.640 ;
        RECT 4.400 302.240 695.600 303.640 ;
        RECT 3.990 300.240 696.000 302.240 ;
        RECT 4.400 298.840 695.600 300.240 ;
        RECT 3.990 296.840 696.000 298.840 ;
        RECT 4.400 295.440 695.600 296.840 ;
        RECT 3.990 293.440 696.000 295.440 ;
        RECT 4.400 292.040 695.600 293.440 ;
        RECT 3.990 290.040 696.000 292.040 ;
        RECT 4.400 288.640 695.600 290.040 ;
        RECT 3.990 286.640 696.000 288.640 ;
        RECT 4.400 285.240 695.600 286.640 ;
        RECT 3.990 283.240 696.000 285.240 ;
        RECT 4.400 281.840 695.600 283.240 ;
        RECT 3.990 279.840 696.000 281.840 ;
        RECT 4.400 278.440 695.600 279.840 ;
        RECT 3.990 276.440 696.000 278.440 ;
        RECT 4.400 275.040 695.600 276.440 ;
        RECT 3.990 273.040 696.000 275.040 ;
        RECT 4.400 271.640 695.600 273.040 ;
        RECT 3.990 269.640 696.000 271.640 ;
        RECT 4.400 268.240 695.600 269.640 ;
        RECT 3.990 266.240 696.000 268.240 ;
        RECT 4.400 264.840 695.600 266.240 ;
        RECT 3.990 262.840 696.000 264.840 ;
        RECT 4.400 261.440 695.600 262.840 ;
        RECT 3.990 259.440 696.000 261.440 ;
        RECT 4.400 258.040 695.600 259.440 ;
        RECT 3.990 256.040 696.000 258.040 ;
        RECT 4.400 254.640 695.600 256.040 ;
        RECT 3.990 252.640 696.000 254.640 ;
        RECT 4.400 251.240 695.600 252.640 ;
        RECT 3.990 249.240 696.000 251.240 ;
        RECT 4.400 247.840 695.600 249.240 ;
        RECT 3.990 245.840 696.000 247.840 ;
        RECT 4.400 244.440 695.600 245.840 ;
        RECT 3.990 242.440 696.000 244.440 ;
        RECT 4.400 241.040 695.600 242.440 ;
        RECT 3.990 239.040 696.000 241.040 ;
        RECT 4.400 237.640 695.600 239.040 ;
        RECT 3.990 235.640 696.000 237.640 ;
        RECT 4.400 234.240 695.600 235.640 ;
        RECT 3.990 232.240 696.000 234.240 ;
        RECT 4.400 230.840 695.600 232.240 ;
        RECT 3.990 228.840 696.000 230.840 ;
        RECT 4.400 227.440 695.600 228.840 ;
        RECT 3.990 225.440 696.000 227.440 ;
        RECT 4.400 224.040 695.600 225.440 ;
        RECT 3.990 222.040 696.000 224.040 ;
        RECT 4.400 220.640 695.600 222.040 ;
        RECT 3.990 218.640 696.000 220.640 ;
        RECT 4.400 217.240 695.600 218.640 ;
        RECT 3.990 215.240 696.000 217.240 ;
        RECT 4.400 213.840 695.600 215.240 ;
        RECT 3.990 211.840 696.000 213.840 ;
        RECT 4.400 210.440 695.600 211.840 ;
        RECT 3.990 208.440 696.000 210.440 ;
        RECT 3.990 207.040 695.600 208.440 ;
        RECT 3.990 205.040 696.000 207.040 ;
        RECT 3.990 203.640 695.600 205.040 ;
        RECT 3.990 201.640 696.000 203.640 ;
        RECT 3.990 200.240 695.600 201.640 ;
        RECT 3.990 198.240 696.000 200.240 ;
        RECT 3.990 196.840 695.600 198.240 ;
        RECT 3.990 194.840 696.000 196.840 ;
        RECT 3.990 193.440 695.600 194.840 ;
        RECT 3.990 191.440 696.000 193.440 ;
        RECT 3.990 190.040 695.600 191.440 ;
        RECT 3.990 188.040 696.000 190.040 ;
        RECT 3.990 186.640 695.600 188.040 ;
        RECT 3.990 184.640 696.000 186.640 ;
        RECT 3.990 183.240 695.600 184.640 ;
        RECT 3.990 181.240 696.000 183.240 ;
        RECT 3.990 179.840 695.600 181.240 ;
        RECT 3.990 177.840 696.000 179.840 ;
        RECT 3.990 176.440 695.600 177.840 ;
        RECT 3.990 174.440 696.000 176.440 ;
        RECT 3.990 173.040 695.600 174.440 ;
        RECT 3.990 171.040 696.000 173.040 ;
        RECT 3.990 169.640 695.600 171.040 ;
        RECT 3.990 167.640 696.000 169.640 ;
        RECT 3.990 166.240 695.600 167.640 ;
        RECT 3.990 164.240 696.000 166.240 ;
        RECT 3.990 162.840 695.600 164.240 ;
        RECT 3.990 160.840 696.000 162.840 ;
        RECT 3.990 159.440 695.600 160.840 ;
        RECT 3.990 157.440 696.000 159.440 ;
        RECT 3.990 156.040 695.600 157.440 ;
        RECT 3.990 154.040 696.000 156.040 ;
        RECT 3.990 152.640 695.600 154.040 ;
        RECT 3.990 150.640 696.000 152.640 ;
        RECT 3.990 149.240 695.600 150.640 ;
        RECT 3.990 147.240 696.000 149.240 ;
        RECT 3.990 145.840 695.600 147.240 ;
        RECT 3.990 143.840 696.000 145.840 ;
        RECT 3.990 142.440 695.600 143.840 ;
        RECT 3.990 140.440 696.000 142.440 ;
        RECT 3.990 139.040 695.600 140.440 ;
        RECT 3.990 137.040 696.000 139.040 ;
        RECT 3.990 135.640 695.600 137.040 ;
        RECT 3.990 133.640 696.000 135.640 ;
        RECT 3.990 132.240 695.600 133.640 ;
        RECT 3.990 130.240 696.000 132.240 ;
        RECT 3.990 128.840 695.600 130.240 ;
        RECT 3.990 126.840 696.000 128.840 ;
        RECT 3.990 125.440 695.600 126.840 ;
        RECT 3.990 123.440 696.000 125.440 ;
        RECT 3.990 122.040 695.600 123.440 ;
        RECT 3.990 120.040 696.000 122.040 ;
        RECT 3.990 118.640 695.600 120.040 ;
        RECT 3.990 116.640 696.000 118.640 ;
        RECT 3.990 115.240 695.600 116.640 ;
        RECT 3.990 113.240 696.000 115.240 ;
        RECT 3.990 111.840 695.600 113.240 ;
        RECT 3.990 109.840 696.000 111.840 ;
        RECT 3.990 108.440 695.600 109.840 ;
        RECT 3.990 106.440 696.000 108.440 ;
        RECT 3.990 105.040 695.600 106.440 ;
        RECT 3.990 103.040 696.000 105.040 ;
        RECT 3.990 101.640 695.600 103.040 ;
        RECT 3.990 99.640 696.000 101.640 ;
        RECT 3.990 98.240 695.600 99.640 ;
        RECT 3.990 96.240 696.000 98.240 ;
        RECT 3.990 94.840 695.600 96.240 ;
        RECT 3.990 35.040 696.000 94.840 ;
        RECT 3.990 33.640 695.600 35.040 ;
        RECT 3.990 10.715 696.000 33.640 ;
      LAYER met4 ;
        RECT 26.975 45.735 174.240 384.705 ;
        RECT 176.640 45.735 177.540 384.705 ;
        RECT 179.940 45.735 327.840 384.705 ;
        RECT 330.240 45.735 331.140 384.705 ;
        RECT 333.540 45.735 481.440 384.705 ;
        RECT 483.840 45.735 484.740 384.705 ;
        RECT 487.140 45.735 635.040 384.705 ;
        RECT 637.440 45.735 638.340 384.705 ;
        RECT 640.740 45.735 679.585 384.705 ;
  END
END team_03
END LIBRARY

